// system_qsys.v

// Generated using ACDS version 13.1 162 at 2019.04.02.17:09:20

`timescale 1 ps / 1 ps
module system_qsys (
		input  wire        clk_clk,                          //                clk.clk
		input  wire        reset_reset_n,                    //              reset.reset_n
		output wire        touch_write,                      //              touch.write
		output wire        touch_read,                       //                   .read
		output wire [31:0] touch_writedata,                  //                   .writedata
		input  wire [31:0] touch_readdata,                   //                   .readdata
		output wire [2:0]  touch_address,                    //                   .address
		output wire        seg_write,                        //                seg.write
		output wire        seg_read,                         //                   .read
		output wire [31:0] seg_writedata,                    //                   .writedata
		input  wire [31:0] seg_readdata,                     //                   .readdata
		output wire [2:0]  seg_address,                      //                   .address
		output wire        remote_write,                     //             remote.write
		output wire        remote_read,                      //                   .read
		output wire [31:0] remote_writedata,                 //                   .writedata
		input  wire [31:0] remote_readdata,                  //                   .readdata
		output wire [2:0]  remote_address,                   //                   .address
		output wire        adda_write,                       //               adda.write
		output wire        adda_read,                        //                   .read
		output wire [31:0] adda_writedata,                   //                   .writedata
		input  wire [31:0] adda_readdata,                    //                   .readdata
		output wire [2:0]  adda_address,                     //                   .address
		input  wire        touch_int_export,                 //          touch_int.export
		input  wire        back_export,                      //               back.export
		input  wire [3:0]  key_export,                       //                key.export
		output wire [3:0]  led_export,                       //                led.export
		output wire        buzzer_export,                    //             buzzer.export
		input  wire        uart_rxd,                         //               uart.rxd
		output wire        uart_txd,                         //                   .txd
		output wire        i2c_scl_export,                   //            i2c_scl.export
		inout  wire        i2c_sda_export,                   //            i2c_sda.export
		input  wire        paint_export,                     //              paint.export
		output wire        ov5640_en_export,                 //          ov5640_en.export
		input  wire        ov5640_id_export,                 //          ov5640_id.export
		output wire        epcs_flash_dclk,                  //         epcs_flash.dclk
		output wire        epcs_flash_sce,                   //                   .sce
		output wire        epcs_flash_sdo,                   //                   .sdo
		input  wire        epcs_flash_data0,                 //                   .data0
		output wire [12:0] sdram_addr,                       //              sdram.addr
		output wire [1:0]  sdram_ba,                         //                   .ba
		output wire        sdram_cas_n,                      //                   .cas_n
		output wire        sdram_cke,                        //                   .cke
		output wire        sdram_cs_n,                       //                   .cs_n
		inout  wire [15:0] sdram_dq,                         //                   .dq
		output wire [1:0]  sdram_dqm,                        //                   .dqm
		output wire        sdram_ras_n,                      //                   .ras_n
		output wire        sdram_we_n,                       //                   .we_n
		output wire        sdram_bridge_slave_waitrequest,   // sdram_bridge_slave.waitrequest
		output wire [15:0] sdram_bridge_slave_readdata,      //                   .readdata
		output wire        sdram_bridge_slave_readdatavalid, //                   .readdatavalid
		input  wire [9:0]  sdram_bridge_slave_burstcount,    //                   .burstcount
		input  wire [15:0] sdram_bridge_slave_writedata,     //                   .writedata
		input  wire [25:0] sdram_bridge_slave_address,       //                   .address
		input  wire        sdram_bridge_slave_write,         //                   .write
		input  wire        sdram_bridge_slave_read,          //                   .read
		input  wire [1:0]  sdram_bridge_slave_byteenable,    //                   .byteenable
		input  wire        sdram_bridge_slave_debugaccess,   //                   .debugaccess
		input  wire [23:0] vip_scl_din_data,                 //        vip_scl_din.data
		input  wire        vip_scl_din_valid,                //                   .valid
		input  wire        vip_scl_din_startofpacket,        //                   .startofpacket
		input  wire        vip_scl_din_endofpacket,          //                   .endofpacket
		output wire        vip_scl_din_ready,                //                   .ready
		output wire [23:0] vip_scl_dout_data,                //       vip_scl_dout.data
		output wire        vip_scl_dout_valid,               //                   .valid
		output wire        vip_scl_dout_startofpacket,       //                   .startofpacket
		output wire        vip_scl_dout_endofpacket,         //                   .endofpacket
		input  wire        vip_scl_dout_ready,               //                   .ready
		output wire        mlcd_cs_n_export,                 //          mlcd_cs_n.export
		output wire        mlcd_wr_n_export,                 //          mlcd_wr_n.export
		output wire        mlcd_rd_n_export,                 //          mlcd_rd_n.export
		output wire        mlcd_rst_n_export,                //         mlcd_rst_n.export
		output wire        mlcd_rs_export,                   //            mlcd_rs.export
		output wire        mlcd_bl_export,                   //            mlcd_bl.export
		input  wire [15:0] lcd_data_in_export,               //        lcd_data_in.export
		output wire [15:0] lcd_data_out_export,              //       lcd_data_out.export
		output wire        lcd_data_dir_export,              //       lcd_data_dir.export
		output wire        lcd_init_done_export,             //      lcd_init_done.export
		output wire [15:0] lcd_id_export,                    //             lcd_id.export
		output wire        eth_mdc_export,                   //            eth_mdc.export
		inout  wire        eth_mdio_export,                  //           eth_mdio.export
		output wire        sd_cs_export,                     //              sd_cs.export
		output wire        sd_clk_export,                    //             sd_clk.export
		output wire        sd_mosi_export,                   //            sd_mosi.export
		input  wire        sd_miso_export,                   //            sd_miso.export
		output wire        page_paint_flag_export,           //    page_paint_flag.export
		output wire        audio_sel_export                  //          audio_sel.export
	);

	wire  [31:0] mm_interconnect_0_pio_page_paint_flag_s1_writedata;        // mm_interconnect_0:pio_page_paint_flag_s1_writedata -> pio_page_paint_flag:writedata
	wire   [1:0] mm_interconnect_0_pio_page_paint_flag_s1_address;          // mm_interconnect_0:pio_page_paint_flag_s1_address -> pio_page_paint_flag:address
	wire         mm_interconnect_0_pio_page_paint_flag_s1_chipselect;       // mm_interconnect_0:pio_page_paint_flag_s1_chipselect -> pio_page_paint_flag:chipselect
	wire         mm_interconnect_0_pio_page_paint_flag_s1_write;            // mm_interconnect_0:pio_page_paint_flag_s1_write -> pio_page_paint_flag:write_n
	wire  [31:0] mm_interconnect_0_pio_page_paint_flag_s1_readdata;         // pio_page_paint_flag:readdata -> mm_interconnect_0:pio_page_paint_flag_s1_readdata
	wire  [31:0] mm_interconnect_0_pio_buzzer_s1_writedata;                 // mm_interconnect_0:pio_buzzer_s1_writedata -> pio_buzzer:writedata
	wire   [1:0] mm_interconnect_0_pio_buzzer_s1_address;                   // mm_interconnect_0:pio_buzzer_s1_address -> pio_buzzer:address
	wire         mm_interconnect_0_pio_buzzer_s1_chipselect;                // mm_interconnect_0:pio_buzzer_s1_chipselect -> pio_buzzer:chipselect
	wire         mm_interconnect_0_pio_buzzer_s1_write;                     // mm_interconnect_0:pio_buzzer_s1_write -> pio_buzzer:write_n
	wire  [31:0] mm_interconnect_0_pio_buzzer_s1_readdata;                  // pio_buzzer:readdata -> mm_interconnect_0:pio_buzzer_s1_readdata
	wire  [31:0] mm_interconnect_0_pio_mlcd_bl_s1_writedata;                // mm_interconnect_0:pio_mlcd_bl_s1_writedata -> pio_mlcd_bl:writedata
	wire   [1:0] mm_interconnect_0_pio_mlcd_bl_s1_address;                  // mm_interconnect_0:pio_mlcd_bl_s1_address -> pio_mlcd_bl:address
	wire         mm_interconnect_0_pio_mlcd_bl_s1_chipselect;               // mm_interconnect_0:pio_mlcd_bl_s1_chipselect -> pio_mlcd_bl:chipselect
	wire         mm_interconnect_0_pio_mlcd_bl_s1_write;                    // mm_interconnect_0:pio_mlcd_bl_s1_write -> pio_mlcd_bl:write_n
	wire  [31:0] mm_interconnect_0_pio_mlcd_bl_s1_readdata;                 // pio_mlcd_bl:readdata -> mm_interconnect_0:pio_mlcd_bl_s1_readdata
	wire  [31:0] mm_interconnect_0_pio_back_s1_writedata;                   // mm_interconnect_0:pio_back_s1_writedata -> pio_back:writedata
	wire   [1:0] mm_interconnect_0_pio_back_s1_address;                     // mm_interconnect_0:pio_back_s1_address -> pio_back:address
	wire         mm_interconnect_0_pio_back_s1_chipselect;                  // mm_interconnect_0:pio_back_s1_chipselect -> pio_back:chipselect
	wire         mm_interconnect_0_pio_back_s1_write;                       // mm_interconnect_0:pio_back_s1_write -> pio_back:write_n
	wire  [31:0] mm_interconnect_0_pio_back_s1_readdata;                    // pio_back:readdata -> mm_interconnect_0:pio_back_s1_readdata
	wire  [31:0] mm_interconnect_0_i2c_scl_s1_writedata;                    // mm_interconnect_0:i2c_scl_s1_writedata -> i2c_scl:writedata
	wire   [1:0] mm_interconnect_0_i2c_scl_s1_address;                      // mm_interconnect_0:i2c_scl_s1_address -> i2c_scl:address
	wire         mm_interconnect_0_i2c_scl_s1_chipselect;                   // mm_interconnect_0:i2c_scl_s1_chipselect -> i2c_scl:chipselect
	wire         mm_interconnect_0_i2c_scl_s1_write;                        // mm_interconnect_0:i2c_scl_s1_write -> i2c_scl:write_n
	wire  [31:0] mm_interconnect_0_i2c_scl_s1_readdata;                     // i2c_scl:readdata -> mm_interconnect_0:i2c_scl_s1_readdata
	wire  [31:0] mm_interconnect_0_pio_mlcd_wr_n_s1_writedata;              // mm_interconnect_0:pio_mlcd_wr_n_s1_writedata -> pio_mlcd_wr_n:writedata
	wire   [1:0] mm_interconnect_0_pio_mlcd_wr_n_s1_address;                // mm_interconnect_0:pio_mlcd_wr_n_s1_address -> pio_mlcd_wr_n:address
	wire         mm_interconnect_0_pio_mlcd_wr_n_s1_chipselect;             // mm_interconnect_0:pio_mlcd_wr_n_s1_chipselect -> pio_mlcd_wr_n:chipselect
	wire         mm_interconnect_0_pio_mlcd_wr_n_s1_write;                  // mm_interconnect_0:pio_mlcd_wr_n_s1_write -> pio_mlcd_wr_n:write_n
	wire  [31:0] mm_interconnect_0_pio_mlcd_wr_n_s1_readdata;               // pio_mlcd_wr_n:readdata -> mm_interconnect_0:pio_mlcd_wr_n_s1_readdata
	wire  [31:0] mm_interconnect_0_pio_lcd_data_out_s1_writedata;           // mm_interconnect_0:pio_lcd_data_out_s1_writedata -> pio_lcd_data_out:writedata
	wire   [1:0] mm_interconnect_0_pio_lcd_data_out_s1_address;             // mm_interconnect_0:pio_lcd_data_out_s1_address -> pio_lcd_data_out:address
	wire         mm_interconnect_0_pio_lcd_data_out_s1_chipselect;          // mm_interconnect_0:pio_lcd_data_out_s1_chipselect -> pio_lcd_data_out:chipselect
	wire         mm_interconnect_0_pio_lcd_data_out_s1_write;               // mm_interconnect_0:pio_lcd_data_out_s1_write -> pio_lcd_data_out:write_n
	wire  [31:0] mm_interconnect_0_pio_lcd_data_out_s1_readdata;            // pio_lcd_data_out:readdata -> mm_interconnect_0:pio_lcd_data_out_s1_readdata
	wire  [31:0] mm_interconnect_0_i2c_sda_s1_writedata;                    // mm_interconnect_0:i2c_sda_s1_writedata -> i2c_sda:writedata
	wire   [1:0] mm_interconnect_0_i2c_sda_s1_address;                      // mm_interconnect_0:i2c_sda_s1_address -> i2c_sda:address
	wire         mm_interconnect_0_i2c_sda_s1_chipselect;                   // mm_interconnect_0:i2c_sda_s1_chipselect -> i2c_sda:chipselect
	wire         mm_interconnect_0_i2c_sda_s1_write;                        // mm_interconnect_0:i2c_sda_s1_write -> i2c_sda:write_n
	wire  [31:0] mm_interconnect_0_i2c_sda_s1_readdata;                     // i2c_sda:readdata -> mm_interconnect_0:i2c_sda_s1_readdata
	wire  [31:0] mm_interconnect_0_pio_lcd_id_s1_writedata;                 // mm_interconnect_0:pio_lcd_id_s1_writedata -> pio_lcd_id:writedata
	wire   [1:0] mm_interconnect_0_pio_lcd_id_s1_address;                   // mm_interconnect_0:pio_lcd_id_s1_address -> pio_lcd_id:address
	wire         mm_interconnect_0_pio_lcd_id_s1_chipselect;                // mm_interconnect_0:pio_lcd_id_s1_chipselect -> pio_lcd_id:chipselect
	wire         mm_interconnect_0_pio_lcd_id_s1_write;                     // mm_interconnect_0:pio_lcd_id_s1_write -> pio_lcd_id:write_n
	wire  [31:0] mm_interconnect_0_pio_lcd_id_s1_readdata;                  // pio_lcd_id:readdata -> mm_interconnect_0:pio_lcd_id_s1_readdata
	wire  [31:0] mm_interconnect_0_pio_sd_mosi_s1_writedata;                // mm_interconnect_0:pio_sd_mosi_s1_writedata -> pio_sd_mosi:writedata
	wire   [1:0] mm_interconnect_0_pio_sd_mosi_s1_address;                  // mm_interconnect_0:pio_sd_mosi_s1_address -> pio_sd_mosi:address
	wire         mm_interconnect_0_pio_sd_mosi_s1_chipselect;               // mm_interconnect_0:pio_sd_mosi_s1_chipselect -> pio_sd_mosi:chipselect
	wire         mm_interconnect_0_pio_sd_mosi_s1_write;                    // mm_interconnect_0:pio_sd_mosi_s1_write -> pio_sd_mosi:write_n
	wire  [31:0] mm_interconnect_0_pio_sd_mosi_s1_readdata;                 // pio_sd_mosi:readdata -> mm_interconnect_0:pio_sd_mosi_s1_readdata
	wire  [31:0] mm_interconnect_0_pio_lcd_data_dir_s1_writedata;           // mm_interconnect_0:pio_lcd_data_dir_s1_writedata -> pio_lcd_data_dir:writedata
	wire   [1:0] mm_interconnect_0_pio_lcd_data_dir_s1_address;             // mm_interconnect_0:pio_lcd_data_dir_s1_address -> pio_lcd_data_dir:address
	wire         mm_interconnect_0_pio_lcd_data_dir_s1_chipselect;          // mm_interconnect_0:pio_lcd_data_dir_s1_chipselect -> pio_lcd_data_dir:chipselect
	wire         mm_interconnect_0_pio_lcd_data_dir_s1_write;               // mm_interconnect_0:pio_lcd_data_dir_s1_write -> pio_lcd_data_dir:write_n
	wire  [31:0] mm_interconnect_0_pio_lcd_data_dir_s1_readdata;            // pio_lcd_data_dir:readdata -> mm_interconnect_0:pio_lcd_data_dir_s1_readdata
	wire         mm_interconnect_0_nios2_jtag_debug_module_waitrequest;     // nios2:jtag_debug_module_waitrequest -> mm_interconnect_0:nios2_jtag_debug_module_waitrequest
	wire  [31:0] mm_interconnect_0_nios2_jtag_debug_module_writedata;       // mm_interconnect_0:nios2_jtag_debug_module_writedata -> nios2:jtag_debug_module_writedata
	wire   [8:0] mm_interconnect_0_nios2_jtag_debug_module_address;         // mm_interconnect_0:nios2_jtag_debug_module_address -> nios2:jtag_debug_module_address
	wire         mm_interconnect_0_nios2_jtag_debug_module_write;           // mm_interconnect_0:nios2_jtag_debug_module_write -> nios2:jtag_debug_module_write
	wire         mm_interconnect_0_nios2_jtag_debug_module_read;            // mm_interconnect_0:nios2_jtag_debug_module_read -> nios2:jtag_debug_module_read
	wire  [31:0] mm_interconnect_0_nios2_jtag_debug_module_readdata;        // nios2:jtag_debug_module_readdata -> mm_interconnect_0:nios2_jtag_debug_module_readdata
	wire         mm_interconnect_0_nios2_jtag_debug_module_debugaccess;     // mm_interconnect_0:nios2_jtag_debug_module_debugaccess -> nios2:jtag_debug_module_debugaccess
	wire   [3:0] mm_interconnect_0_nios2_jtag_debug_module_byteenable;      // mm_interconnect_0:nios2_jtag_debug_module_byteenable -> nios2:jtag_debug_module_byteenable
	wire  [31:0] mm_interconnect_0_pio_ov5640_en_s1_writedata;              // mm_interconnect_0:pio_ov5640_en_s1_writedata -> pio_ov5640_en:writedata
	wire   [1:0] mm_interconnect_0_pio_ov5640_en_s1_address;                // mm_interconnect_0:pio_ov5640_en_s1_address -> pio_ov5640_en:address
	wire         mm_interconnect_0_pio_ov5640_en_s1_chipselect;             // mm_interconnect_0:pio_ov5640_en_s1_chipselect -> pio_ov5640_en:chipselect
	wire         mm_interconnect_0_pio_ov5640_en_s1_write;                  // mm_interconnect_0:pio_ov5640_en_s1_write -> pio_ov5640_en:write_n
	wire  [31:0] mm_interconnect_0_pio_ov5640_en_s1_readdata;               // pio_ov5640_en:readdata -> mm_interconnect_0:pio_ov5640_en_s1_readdata
	wire  [31:0] mm_interconnect_0_pio_lcd_init_done_s1_writedata;          // mm_interconnect_0:pio_lcd_init_done_s1_writedata -> pio_lcd_init_done:writedata
	wire   [1:0] mm_interconnect_0_pio_lcd_init_done_s1_address;            // mm_interconnect_0:pio_lcd_init_done_s1_address -> pio_lcd_init_done:address
	wire         mm_interconnect_0_pio_lcd_init_done_s1_chipselect;         // mm_interconnect_0:pio_lcd_init_done_s1_chipselect -> pio_lcd_init_done:chipselect
	wire         mm_interconnect_0_pio_lcd_init_done_s1_write;              // mm_interconnect_0:pio_lcd_init_done_s1_write -> pio_lcd_init_done:write_n
	wire  [31:0] mm_interconnect_0_pio_lcd_init_done_s1_readdata;           // pio_lcd_init_done:readdata -> mm_interconnect_0:pio_lcd_init_done_s1_readdata
	wire   [1:0] mm_interconnect_0_pio_ov5640_id_s1_address;                // mm_interconnect_0:pio_ov5640_id_s1_address -> pio_ov5640_id:address
	wire  [31:0] mm_interconnect_0_pio_ov5640_id_s1_readdata;               // pio_ov5640_id:readdata -> mm_interconnect_0:pio_ov5640_id_s1_readdata
	wire         nios2_data_master_waitrequest;                             // mm_interconnect_0:nios2_data_master_waitrequest -> nios2:d_waitrequest
	wire  [31:0] nios2_data_master_writedata;                               // nios2:d_writedata -> mm_interconnect_0:nios2_data_master_writedata
	wire  [25:0] nios2_data_master_address;                                 // nios2:d_address -> mm_interconnect_0:nios2_data_master_address
	wire         nios2_data_master_write;                                   // nios2:d_write -> mm_interconnect_0:nios2_data_master_write
	wire         nios2_data_master_read;                                    // nios2:d_read -> mm_interconnect_0:nios2_data_master_read
	wire  [31:0] nios2_data_master_readdata;                                // mm_interconnect_0:nios2_data_master_readdata -> nios2:d_readdata
	wire         nios2_data_master_debugaccess;                             // nios2:jtag_debug_module_debugaccess_to_roms -> mm_interconnect_0:nios2_data_master_debugaccess
	wire         nios2_data_master_readdatavalid;                           // mm_interconnect_0:nios2_data_master_readdatavalid -> nios2:d_readdatavalid
	wire   [3:0] nios2_data_master_byteenable;                              // nios2:d_byteenable -> mm_interconnect_0:nios2_data_master_byteenable
	wire   [9:0] sdram_bridge_m0_burstcount;                                // sdram_bridge:m0_burstcount -> mm_interconnect_0:sdram_bridge_m0_burstcount
	wire         sdram_bridge_m0_waitrequest;                               // mm_interconnect_0:sdram_bridge_m0_waitrequest -> sdram_bridge:m0_waitrequest
	wire  [25:0] sdram_bridge_m0_address;                                   // sdram_bridge:m0_address -> mm_interconnect_0:sdram_bridge_m0_address
	wire  [15:0] sdram_bridge_m0_writedata;                                 // sdram_bridge:m0_writedata -> mm_interconnect_0:sdram_bridge_m0_writedata
	wire         sdram_bridge_m0_write;                                     // sdram_bridge:m0_write -> mm_interconnect_0:sdram_bridge_m0_write
	wire         sdram_bridge_m0_read;                                      // sdram_bridge:m0_read -> mm_interconnect_0:sdram_bridge_m0_read
	wire  [15:0] sdram_bridge_m0_readdata;                                  // mm_interconnect_0:sdram_bridge_m0_readdata -> sdram_bridge:m0_readdata
	wire         sdram_bridge_m0_debugaccess;                               // sdram_bridge:m0_debugaccess -> mm_interconnect_0:sdram_bridge_m0_debugaccess
	wire   [1:0] sdram_bridge_m0_byteenable;                                // sdram_bridge:m0_byteenable -> mm_interconnect_0:sdram_bridge_m0_byteenable
	wire         sdram_bridge_m0_readdatavalid;                             // mm_interconnect_0:sdram_bridge_m0_readdatavalid -> sdram_bridge:m0_readdatavalid
	wire  [31:0] mm_interconnect_0_mm_bridge_adda_avalon_slave_writedata;   // mm_interconnect_0:mm_bridge_adda_avalon_slave_writedata -> mm_bridge_adda:avalon_writedata
	wire   [2:0] mm_interconnect_0_mm_bridge_adda_avalon_slave_address;     // mm_interconnect_0:mm_bridge_adda_avalon_slave_address -> mm_bridge_adda:avalon_address
	wire         mm_interconnect_0_mm_bridge_adda_avalon_slave_write;       // mm_interconnect_0:mm_bridge_adda_avalon_slave_write -> mm_bridge_adda:avalon_write
	wire         mm_interconnect_0_mm_bridge_adda_avalon_slave_read;        // mm_interconnect_0:mm_bridge_adda_avalon_slave_read -> mm_bridge_adda:avalon_read
	wire  [31:0] mm_interconnect_0_mm_bridge_adda_avalon_slave_readdata;    // mm_bridge_adda:avalon_readdata -> mm_interconnect_0:mm_bridge_adda_avalon_slave_readdata
	wire  [31:0] mm_interconnect_0_pio_touch_int_s1_writedata;              // mm_interconnect_0:pio_touch_int_s1_writedata -> pio_touch_int:writedata
	wire   [1:0] mm_interconnect_0_pio_touch_int_s1_address;                // mm_interconnect_0:pio_touch_int_s1_address -> pio_touch_int:address
	wire         mm_interconnect_0_pio_touch_int_s1_chipselect;             // mm_interconnect_0:pio_touch_int_s1_chipselect -> pio_touch_int:chipselect
	wire         mm_interconnect_0_pio_touch_int_s1_write;                  // mm_interconnect_0:pio_touch_int_s1_write -> pio_touch_int:write_n
	wire  [31:0] mm_interconnect_0_pio_touch_int_s1_readdata;               // pio_touch_int:readdata -> mm_interconnect_0:pio_touch_int_s1_readdata
	wire  [31:0] mm_interconnect_0_pio_mlcd_cs_n_s1_writedata;              // mm_interconnect_0:pio_mlcd_cs_n_s1_writedata -> pio_mlcd_cs_n:writedata
	wire   [1:0] mm_interconnect_0_pio_mlcd_cs_n_s1_address;                // mm_interconnect_0:pio_mlcd_cs_n_s1_address -> pio_mlcd_cs_n:address
	wire         mm_interconnect_0_pio_mlcd_cs_n_s1_chipselect;             // mm_interconnect_0:pio_mlcd_cs_n_s1_chipselect -> pio_mlcd_cs_n:chipselect
	wire         mm_interconnect_0_pio_mlcd_cs_n_s1_write;                  // mm_interconnect_0:pio_mlcd_cs_n_s1_write -> pio_mlcd_cs_n:write_n
	wire  [31:0] mm_interconnect_0_pio_mlcd_cs_n_s1_readdata;               // pio_mlcd_cs_n:readdata -> mm_interconnect_0:pio_mlcd_cs_n_s1_readdata
	wire  [31:0] mm_interconnect_0_mm_bridge_touch_avalon_slave_writedata;  // mm_interconnect_0:mm_bridge_touch_avalon_slave_writedata -> mm_bridge_touch:avalon_writedata
	wire   [2:0] mm_interconnect_0_mm_bridge_touch_avalon_slave_address;    // mm_interconnect_0:mm_bridge_touch_avalon_slave_address -> mm_bridge_touch:avalon_address
	wire         mm_interconnect_0_mm_bridge_touch_avalon_slave_write;      // mm_interconnect_0:mm_bridge_touch_avalon_slave_write -> mm_bridge_touch:avalon_write
	wire         mm_interconnect_0_mm_bridge_touch_avalon_slave_read;       // mm_interconnect_0:mm_bridge_touch_avalon_slave_read -> mm_bridge_touch:avalon_read
	wire  [31:0] mm_interconnect_0_mm_bridge_touch_avalon_slave_readdata;   // mm_bridge_touch:avalon_readdata -> mm_interconnect_0:mm_bridge_touch_avalon_slave_readdata
	wire   [0:0] mm_interconnect_0_sysid_control_slave_address;             // mm_interconnect_0:sysid_control_slave_address -> sysid:address
	wire  [31:0] mm_interconnect_0_sysid_control_slave_readdata;            // sysid:readdata -> mm_interconnect_0:sysid_control_slave_readdata
	wire  [31:0] mm_interconnect_0_pio_mdc_s1_writedata;                    // mm_interconnect_0:pio_mdc_s1_writedata -> pio_mdc:writedata
	wire   [1:0] mm_interconnect_0_pio_mdc_s1_address;                      // mm_interconnect_0:pio_mdc_s1_address -> pio_mdc:address
	wire         mm_interconnect_0_pio_mdc_s1_chipselect;                   // mm_interconnect_0:pio_mdc_s1_chipselect -> pio_mdc:chipselect
	wire         mm_interconnect_0_pio_mdc_s1_write;                        // mm_interconnect_0:pio_mdc_s1_write -> pio_mdc:write_n
	wire  [31:0] mm_interconnect_0_pio_mdc_s1_readdata;                     // pio_mdc:readdata -> mm_interconnect_0:pio_mdc_s1_readdata
	wire  [31:0] mm_interconnect_0_pio_mlcd_rd_n_s1_writedata;              // mm_interconnect_0:pio_mlcd_rd_n_s1_writedata -> pio_mlcd_rd_n:writedata
	wire   [1:0] mm_interconnect_0_pio_mlcd_rd_n_s1_address;                // mm_interconnect_0:pio_mlcd_rd_n_s1_address -> pio_mlcd_rd_n:address
	wire         mm_interconnect_0_pio_mlcd_rd_n_s1_chipselect;             // mm_interconnect_0:pio_mlcd_rd_n_s1_chipselect -> pio_mlcd_rd_n:chipselect
	wire         mm_interconnect_0_pio_mlcd_rd_n_s1_write;                  // mm_interconnect_0:pio_mlcd_rd_n_s1_write -> pio_mlcd_rd_n:write_n
	wire  [31:0] mm_interconnect_0_pio_mlcd_rd_n_s1_readdata;               // pio_mlcd_rd_n:readdata -> mm_interconnect_0:pio_mlcd_rd_n_s1_readdata
	wire  [31:0] mm_interconnect_0_pio_mdio_s1_writedata;                   // mm_interconnect_0:pio_mdio_s1_writedata -> pio_mdio:writedata
	wire   [1:0] mm_interconnect_0_pio_mdio_s1_address;                     // mm_interconnect_0:pio_mdio_s1_address -> pio_mdio:address
	wire         mm_interconnect_0_pio_mdio_s1_chipselect;                  // mm_interconnect_0:pio_mdio_s1_chipselect -> pio_mdio:chipselect
	wire         mm_interconnect_0_pio_mdio_s1_write;                       // mm_interconnect_0:pio_mdio_s1_write -> pio_mdio:write_n
	wire  [31:0] mm_interconnect_0_pio_mdio_s1_readdata;                    // pio_mdio:readdata -> mm_interconnect_0:pio_mdio_s1_readdata
	wire         nios2_instruction_master_waitrequest;                      // mm_interconnect_0:nios2_instruction_master_waitrequest -> nios2:i_waitrequest
	wire  [25:0] nios2_instruction_master_address;                          // nios2:i_address -> mm_interconnect_0:nios2_instruction_master_address
	wire         nios2_instruction_master_read;                             // nios2:i_read -> mm_interconnect_0:nios2_instruction_master_read
	wire  [31:0] nios2_instruction_master_readdata;                         // mm_interconnect_0:nios2_instruction_master_readdata -> nios2:i_readdata
	wire         nios2_instruction_master_readdatavalid;                    // mm_interconnect_0:nios2_instruction_master_readdatavalid -> nios2:i_readdatavalid
	wire  [31:0] mm_interconnect_0_mm_bridge_seg_avalon_slave_writedata;    // mm_interconnect_0:mm_bridge_seg_avalon_slave_writedata -> mm_bridge_seg:avalon_writedata
	wire   [2:0] mm_interconnect_0_mm_bridge_seg_avalon_slave_address;      // mm_interconnect_0:mm_bridge_seg_avalon_slave_address -> mm_bridge_seg:avalon_address
	wire         mm_interconnect_0_mm_bridge_seg_avalon_slave_write;        // mm_interconnect_0:mm_bridge_seg_avalon_slave_write -> mm_bridge_seg:avalon_write
	wire         mm_interconnect_0_mm_bridge_seg_avalon_slave_read;         // mm_interconnect_0:mm_bridge_seg_avalon_slave_read -> mm_bridge_seg:avalon_read
	wire  [31:0] mm_interconnect_0_mm_bridge_seg_avalon_slave_readdata;     // mm_bridge_seg:avalon_readdata -> mm_interconnect_0:mm_bridge_seg_avalon_slave_readdata
	wire         mm_interconnect_0_alt_vip_cl_scl_0_control_waitrequest;    // alt_vip_cl_scl_0:control_waitrequest -> mm_interconnect_0:alt_vip_cl_scl_0_control_waitrequest
	wire  [31:0] mm_interconnect_0_alt_vip_cl_scl_0_control_writedata;      // mm_interconnect_0:alt_vip_cl_scl_0_control_writedata -> alt_vip_cl_scl_0:control_writedata
	wire   [6:0] mm_interconnect_0_alt_vip_cl_scl_0_control_address;        // mm_interconnect_0:alt_vip_cl_scl_0_control_address -> alt_vip_cl_scl_0:control_address
	wire         mm_interconnect_0_alt_vip_cl_scl_0_control_write;          // mm_interconnect_0:alt_vip_cl_scl_0_control_write -> alt_vip_cl_scl_0:control_write
	wire         mm_interconnect_0_alt_vip_cl_scl_0_control_read;           // mm_interconnect_0:alt_vip_cl_scl_0_control_read -> alt_vip_cl_scl_0:control_read
	wire  [31:0] mm_interconnect_0_alt_vip_cl_scl_0_control_readdata;       // alt_vip_cl_scl_0:control_readdata -> mm_interconnect_0:alt_vip_cl_scl_0_control_readdata
	wire         mm_interconnect_0_alt_vip_cl_scl_0_control_readdatavalid;  // alt_vip_cl_scl_0:control_readdatavalid -> mm_interconnect_0:alt_vip_cl_scl_0_control_readdatavalid
	wire   [3:0] mm_interconnect_0_alt_vip_cl_scl_0_control_byteenable;     // mm_interconnect_0:alt_vip_cl_scl_0_control_byteenable -> alt_vip_cl_scl_0:control_byteenable
	wire  [31:0] mm_interconnect_0_pio_sd_clk_s1_writedata;                 // mm_interconnect_0:pio_sd_clk_s1_writedata -> pio_sd_clk:writedata
	wire   [1:0] mm_interconnect_0_pio_sd_clk_s1_address;                   // mm_interconnect_0:pio_sd_clk_s1_address -> pio_sd_clk:address
	wire         mm_interconnect_0_pio_sd_clk_s1_chipselect;                // mm_interconnect_0:pio_sd_clk_s1_chipselect -> pio_sd_clk:chipselect
	wire         mm_interconnect_0_pio_sd_clk_s1_write;                     // mm_interconnect_0:pio_sd_clk_s1_write -> pio_sd_clk:write_n
	wire  [31:0] mm_interconnect_0_pio_sd_clk_s1_readdata;                  // pio_sd_clk:readdata -> mm_interconnect_0:pio_sd_clk_s1_readdata
	wire  [31:0] mm_interconnect_0_pio_mlcd_rst_n_s1_writedata;             // mm_interconnect_0:pio_mlcd_rst_n_s1_writedata -> pio_mlcd_rst_n:writedata
	wire   [1:0] mm_interconnect_0_pio_mlcd_rst_n_s1_address;               // mm_interconnect_0:pio_mlcd_rst_n_s1_address -> pio_mlcd_rst_n:address
	wire         mm_interconnect_0_pio_mlcd_rst_n_s1_chipselect;            // mm_interconnect_0:pio_mlcd_rst_n_s1_chipselect -> pio_mlcd_rst_n:chipselect
	wire         mm_interconnect_0_pio_mlcd_rst_n_s1_write;                 // mm_interconnect_0:pio_mlcd_rst_n_s1_write -> pio_mlcd_rst_n:write_n
	wire  [31:0] mm_interconnect_0_pio_mlcd_rst_n_s1_readdata;              // pio_mlcd_rst_n:readdata -> mm_interconnect_0:pio_mlcd_rst_n_s1_readdata
	wire  [31:0] mm_interconnect_0_pio_paint_s1_writedata;                  // mm_interconnect_0:pio_paint_s1_writedata -> pio_paint:writedata
	wire   [1:0] mm_interconnect_0_pio_paint_s1_address;                    // mm_interconnect_0:pio_paint_s1_address -> pio_paint:address
	wire         mm_interconnect_0_pio_paint_s1_chipselect;                 // mm_interconnect_0:pio_paint_s1_chipselect -> pio_paint:chipselect
	wire         mm_interconnect_0_pio_paint_s1_write;                      // mm_interconnect_0:pio_paint_s1_write -> pio_paint:write_n
	wire  [31:0] mm_interconnect_0_pio_paint_s1_readdata;                   // pio_paint:readdata -> mm_interconnect_0:pio_paint_s1_readdata
	wire   [1:0] mm_interconnect_0_pio_lcd_data_in_s1_address;              // mm_interconnect_0:pio_lcd_data_in_s1_address -> pio_lcd_data_in:address
	wire  [31:0] mm_interconnect_0_pio_lcd_data_in_s1_readdata;             // pio_lcd_data_in:readdata -> mm_interconnect_0:pio_lcd_data_in_s1_readdata
	wire   [1:0] mm_interconnect_0_pio_key_s1_address;                      // mm_interconnect_0:pio_key_s1_address -> pio_key:address
	wire  [31:0] mm_interconnect_0_pio_key_s1_readdata;                     // pio_key:readdata -> mm_interconnect_0:pio_key_s1_readdata
	wire  [31:0] mm_interconnect_0_pio_sd_cs_s1_writedata;                  // mm_interconnect_0:pio_sd_cs_s1_writedata -> pio_sd_cs:writedata
	wire   [1:0] mm_interconnect_0_pio_sd_cs_s1_address;                    // mm_interconnect_0:pio_sd_cs_s1_address -> pio_sd_cs:address
	wire         mm_interconnect_0_pio_sd_cs_s1_chipselect;                 // mm_interconnect_0:pio_sd_cs_s1_chipselect -> pio_sd_cs:chipselect
	wire         mm_interconnect_0_pio_sd_cs_s1_write;                      // mm_interconnect_0:pio_sd_cs_s1_write -> pio_sd_cs:write_n
	wire  [31:0] mm_interconnect_0_pio_sd_cs_s1_readdata;                   // pio_sd_cs:readdata -> mm_interconnect_0:pio_sd_cs_s1_readdata
	wire  [31:0] mm_interconnect_0_pio_led_s1_writedata;                    // mm_interconnect_0:pio_led_s1_writedata -> pio_led:writedata
	wire   [1:0] mm_interconnect_0_pio_led_s1_address;                      // mm_interconnect_0:pio_led_s1_address -> pio_led:address
	wire         mm_interconnect_0_pio_led_s1_chipselect;                   // mm_interconnect_0:pio_led_s1_chipselect -> pio_led:chipselect
	wire         mm_interconnect_0_pio_led_s1_write;                        // mm_interconnect_0:pio_led_s1_write -> pio_led:write_n
	wire  [31:0] mm_interconnect_0_pio_led_s1_readdata;                     // pio_led:readdata -> mm_interconnect_0:pio_led_s1_readdata
	wire   [1:0] mm_interconnect_0_pio_sd_miso_s1_address;                  // mm_interconnect_0:pio_sd_miso_s1_address -> pio_sd_miso:address
	wire  [31:0] mm_interconnect_0_pio_sd_miso_s1_readdata;                 // pio_sd_miso:readdata -> mm_interconnect_0:pio_sd_miso_s1_readdata
	wire         mm_interconnect_0_sdram_s1_waitrequest;                    // sdram:za_waitrequest -> mm_interconnect_0:sdram_s1_waitrequest
	wire  [15:0] mm_interconnect_0_sdram_s1_writedata;                      // mm_interconnect_0:sdram_s1_writedata -> sdram:az_data
	wire  [23:0] mm_interconnect_0_sdram_s1_address;                        // mm_interconnect_0:sdram_s1_address -> sdram:az_addr
	wire         mm_interconnect_0_sdram_s1_chipselect;                     // mm_interconnect_0:sdram_s1_chipselect -> sdram:az_cs
	wire         mm_interconnect_0_sdram_s1_write;                          // mm_interconnect_0:sdram_s1_write -> sdram:az_wr_n
	wire         mm_interconnect_0_sdram_s1_read;                           // mm_interconnect_0:sdram_s1_read -> sdram:az_rd_n
	wire  [15:0] mm_interconnect_0_sdram_s1_readdata;                       // sdram:za_data -> mm_interconnect_0:sdram_s1_readdata
	wire         mm_interconnect_0_sdram_s1_readdatavalid;                  // sdram:za_valid -> mm_interconnect_0:sdram_s1_readdatavalid
	wire   [1:0] mm_interconnect_0_sdram_s1_byteenable;                     // mm_interconnect_0:sdram_s1_byteenable -> sdram:az_be_n
	wire  [31:0] mm_interconnect_0_pio_mlcd_rs_s1_writedata;                // mm_interconnect_0:pio_mlcd_rs_s1_writedata -> pio_mlcd_rs:writedata
	wire   [1:0] mm_interconnect_0_pio_mlcd_rs_s1_address;                  // mm_interconnect_0:pio_mlcd_rs_s1_address -> pio_mlcd_rs:address
	wire         mm_interconnect_0_pio_mlcd_rs_s1_chipselect;               // mm_interconnect_0:pio_mlcd_rs_s1_chipselect -> pio_mlcd_rs:chipselect
	wire         mm_interconnect_0_pio_mlcd_rs_s1_write;                    // mm_interconnect_0:pio_mlcd_rs_s1_write -> pio_mlcd_rs:write_n
	wire  [31:0] mm_interconnect_0_pio_mlcd_rs_s1_readdata;                 // pio_mlcd_rs:readdata -> mm_interconnect_0:pio_mlcd_rs_s1_readdata
	wire  [31:0] mm_interconnect_0_pio_audio_sel_s1_writedata;              // mm_interconnect_0:pio_audio_sel_s1_writedata -> pio_audio_sel:writedata
	wire   [1:0] mm_interconnect_0_pio_audio_sel_s1_address;                // mm_interconnect_0:pio_audio_sel_s1_address -> pio_audio_sel:address
	wire         mm_interconnect_0_pio_audio_sel_s1_chipselect;             // mm_interconnect_0:pio_audio_sel_s1_chipselect -> pio_audio_sel:chipselect
	wire         mm_interconnect_0_pio_audio_sel_s1_write;                  // mm_interconnect_0:pio_audio_sel_s1_write -> pio_audio_sel:write_n
	wire  [31:0] mm_interconnect_0_pio_audio_sel_s1_readdata;               // pio_audio_sel:readdata -> mm_interconnect_0:pio_audio_sel_s1_readdata
	wire  [31:0] mm_interconnect_0_mm_bridge_remote_avalon_slave_writedata; // mm_interconnect_0:mm_bridge_remote_avalon_slave_writedata -> mm_bridge_remote:avalon_writedata
	wire   [2:0] mm_interconnect_0_mm_bridge_remote_avalon_slave_address;   // mm_interconnect_0:mm_bridge_remote_avalon_slave_address -> mm_bridge_remote:avalon_address
	wire         mm_interconnect_0_mm_bridge_remote_avalon_slave_write;     // mm_interconnect_0:mm_bridge_remote_avalon_slave_write -> mm_bridge_remote:avalon_write
	wire         mm_interconnect_0_mm_bridge_remote_avalon_slave_read;      // mm_interconnect_0:mm_bridge_remote_avalon_slave_read -> mm_bridge_remote:avalon_read
	wire  [31:0] mm_interconnect_0_mm_bridge_remote_avalon_slave_readdata;  // mm_bridge_remote:avalon_readdata -> mm_interconnect_0:mm_bridge_remote_avalon_slave_readdata
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest; // jtag_uart:av_waitrequest -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_waitrequest
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata;   // mm_interconnect_0:jtag_uart_avalon_jtag_slave_writedata -> jtag_uart:av_writedata
	wire   [0:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_address;     // mm_interconnect_0:jtag_uart_avalon_jtag_slave_address -> jtag_uart:av_address
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect;  // mm_interconnect_0:jtag_uart_avalon_jtag_slave_chipselect -> jtag_uart:av_chipselect
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_write;       // mm_interconnect_0:jtag_uart_avalon_jtag_slave_write -> jtag_uart:av_write_n
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_read;        // mm_interconnect_0:jtag_uart_avalon_jtag_slave_read -> jtag_uart:av_read_n
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata;    // jtag_uart:av_readdata -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_readdata
	wire  [31:0] mm_interconnect_0_epcs_flash_epcs_control_port_writedata;  // mm_interconnect_0:epcs_flash_epcs_control_port_writedata -> epcs_flash:writedata
	wire   [8:0] mm_interconnect_0_epcs_flash_epcs_control_port_address;    // mm_interconnect_0:epcs_flash_epcs_control_port_address -> epcs_flash:address
	wire         mm_interconnect_0_epcs_flash_epcs_control_port_chipselect; // mm_interconnect_0:epcs_flash_epcs_control_port_chipselect -> epcs_flash:chipselect
	wire         mm_interconnect_0_epcs_flash_epcs_control_port_write;      // mm_interconnect_0:epcs_flash_epcs_control_port_write -> epcs_flash:write_n
	wire         mm_interconnect_0_epcs_flash_epcs_control_port_read;       // mm_interconnect_0:epcs_flash_epcs_control_port_read -> epcs_flash:read_n
	wire  [31:0] mm_interconnect_0_epcs_flash_epcs_control_port_readdata;   // epcs_flash:readdata -> mm_interconnect_0:epcs_flash_epcs_control_port_readdata
	wire  [15:0] mm_interconnect_0_uart_s1_writedata;                       // mm_interconnect_0:uart_s1_writedata -> uart:writedata
	wire   [2:0] mm_interconnect_0_uart_s1_address;                         // mm_interconnect_0:uart_s1_address -> uart:address
	wire         mm_interconnect_0_uart_s1_chipselect;                      // mm_interconnect_0:uart_s1_chipselect -> uart:chipselect
	wire         mm_interconnect_0_uart_s1_write;                           // mm_interconnect_0:uart_s1_write -> uart:write_n
	wire         mm_interconnect_0_uart_s1_read;                            // mm_interconnect_0:uart_s1_read -> uart:read_n
	wire  [15:0] mm_interconnect_0_uart_s1_readdata;                        // uart:readdata -> mm_interconnect_0:uart_s1_readdata
	wire         mm_interconnect_0_uart_s1_begintransfer;                   // mm_interconnect_0:uart_s1_begintransfer -> uart:begintransfer
	wire         irq_mapper_receiver0_irq;                                  // jtag_uart:av_irq -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                                  // epcs_flash:irq -> irq_mapper:receiver1_irq
	wire         irq_mapper_receiver2_irq;                                  // uart:irq -> irq_mapper:receiver2_irq
	wire         irq_mapper_receiver3_irq;                                  // pio_touch_int:irq -> irq_mapper:receiver3_irq
	wire         irq_mapper_receiver4_irq;                                  // pio_back:irq -> irq_mapper:receiver4_irq
	wire         irq_mapper_receiver5_irq;                                  // pio_paint:irq -> irq_mapper:receiver5_irq
	wire  [31:0] nios2_d_irq_irq;                                           // irq_mapper:sender_irq -> nios2:d_irq
	wire         rst_controller_reset_out_reset;                            // rst_controller:reset_out -> [alt_vip_cl_scl_0:main_reset, epcs_flash:reset_n, i2c_scl:reset_n, i2c_sda:reset_n, irq_mapper:reset, jtag_uart:rst_n, mm_bridge_adda:rst_n, mm_bridge_remote:rst_n, mm_bridge_seg:rst_n, mm_bridge_touch:rst_n, mm_interconnect_0:nios2_reset_n_reset_bridge_in_reset_reset, nios2:reset_n, pio_audio_sel:reset_n, pio_back:reset_n, pio_buzzer:reset_n, pio_key:reset_n, pio_lcd_data_dir:reset_n, pio_lcd_data_in:reset_n, pio_lcd_data_out:reset_n, pio_lcd_id:reset_n, pio_lcd_init_done:reset_n, pio_led:reset_n, pio_mdc:reset_n, pio_mdio:reset_n, pio_mlcd_bl:reset_n, pio_mlcd_cs_n:reset_n, pio_mlcd_rd_n:reset_n, pio_mlcd_rs:reset_n, pio_mlcd_rst_n:reset_n, pio_mlcd_wr_n:reset_n, pio_ov5640_en:reset_n, pio_ov5640_id:reset_n, pio_page_paint_flag:reset_n, pio_paint:reset_n, pio_sd_clk:reset_n, pio_sd_cs:reset_n, pio_sd_miso:reset_n, pio_sd_mosi:reset_n, pio_touch_int:reset_n, rst_translator:in_reset, sdram:reset_n, sdram_bridge:reset, sysid:reset_n, uart:reset_n]
	wire         rst_controller_reset_out_reset_req;                        // rst_controller:reset_req -> [epcs_flash:reset_req, nios2:reset_req, rst_translator:reset_req_in]
	wire         nios2_jtag_debug_module_reset_reset;                       // nios2:jtag_debug_module_resetrequest -> rst_controller:reset_in1

	system_qsys_nios2 nios2 (
		.clk                                   (clk_clk),                                               //                       clk.clk
		.reset_n                               (~rst_controller_reset_out_reset),                       //                   reset_n.reset_n
		.reset_req                             (rst_controller_reset_out_reset_req),                    //                          .reset_req
		.d_address                             (nios2_data_master_address),                             //               data_master.address
		.d_byteenable                          (nios2_data_master_byteenable),                          //                          .byteenable
		.d_read                                (nios2_data_master_read),                                //                          .read
		.d_readdata                            (nios2_data_master_readdata),                            //                          .readdata
		.d_waitrequest                         (nios2_data_master_waitrequest),                         //                          .waitrequest
		.d_write                               (nios2_data_master_write),                               //                          .write
		.d_writedata                           (nios2_data_master_writedata),                           //                          .writedata
		.d_readdatavalid                       (nios2_data_master_readdatavalid),                       //                          .readdatavalid
		.jtag_debug_module_debugaccess_to_roms (nios2_data_master_debugaccess),                         //                          .debugaccess
		.i_address                             (nios2_instruction_master_address),                      //        instruction_master.address
		.i_read                                (nios2_instruction_master_read),                         //                          .read
		.i_readdata                            (nios2_instruction_master_readdata),                     //                          .readdata
		.i_waitrequest                         (nios2_instruction_master_waitrequest),                  //                          .waitrequest
		.i_readdatavalid                       (nios2_instruction_master_readdatavalid),                //                          .readdatavalid
		.d_irq                                 (nios2_d_irq_irq),                                       //                     d_irq.irq
		.jtag_debug_module_resetrequest        (nios2_jtag_debug_module_reset_reset),                   //   jtag_debug_module_reset.reset
		.jtag_debug_module_address             (mm_interconnect_0_nios2_jtag_debug_module_address),     //         jtag_debug_module.address
		.jtag_debug_module_byteenable          (mm_interconnect_0_nios2_jtag_debug_module_byteenable),  //                          .byteenable
		.jtag_debug_module_debugaccess         (mm_interconnect_0_nios2_jtag_debug_module_debugaccess), //                          .debugaccess
		.jtag_debug_module_read                (mm_interconnect_0_nios2_jtag_debug_module_read),        //                          .read
		.jtag_debug_module_readdata            (mm_interconnect_0_nios2_jtag_debug_module_readdata),    //                          .readdata
		.jtag_debug_module_waitrequest         (mm_interconnect_0_nios2_jtag_debug_module_waitrequest), //                          .waitrequest
		.jtag_debug_module_write               (mm_interconnect_0_nios2_jtag_debug_module_write),       //                          .write
		.jtag_debug_module_writedata           (mm_interconnect_0_nios2_jtag_debug_module_writedata),   //                          .writedata
		.no_ci_readra                          ()                                                       // custom_instruction_master.readra
	);

	system_qsys_jtag_uart jtag_uart (
		.clk            (clk_clk),                                                   //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                           //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver0_irq)                                   //               irq.irq
	);

	system_qsys_epcs_flash epcs_flash (
		.clk           (clk_clk),                                                   //               clk.clk
		.reset_n       (~rst_controller_reset_out_reset),                           //             reset.reset_n
		.reset_req     (rst_controller_reset_out_reset_req),                        //                  .reset_req
		.address       (mm_interconnect_0_epcs_flash_epcs_control_port_address),    // epcs_control_port.address
		.chipselect    (mm_interconnect_0_epcs_flash_epcs_control_port_chipselect), //                  .chipselect
		.dataavailable (),                                                          //                  .dataavailable
		.endofpacket   (),                                                          //                  .endofpacket
		.read_n        (~mm_interconnect_0_epcs_flash_epcs_control_port_read),      //                  .read_n
		.readdata      (mm_interconnect_0_epcs_flash_epcs_control_port_readdata),   //                  .readdata
		.readyfordata  (),                                                          //                  .readyfordata
		.write_n       (~mm_interconnect_0_epcs_flash_epcs_control_port_write),     //                  .write_n
		.writedata     (mm_interconnect_0_epcs_flash_epcs_control_port_writedata),  //                  .writedata
		.irq           (irq_mapper_receiver1_irq),                                  //               irq.irq
		.dclk          (epcs_flash_dclk),                                           //          external.export
		.sce           (epcs_flash_sce),                                            //                  .export
		.sdo           (epcs_flash_sdo),                                            //                  .export
		.data0         (epcs_flash_data0)                                           //                  .export
	);

	system_qsys_sdram sdram (
		.clk            (clk_clk),                                  //   clk.clk
		.reset_n        (~rst_controller_reset_out_reset),          // reset.reset_n
		.az_addr        (mm_interconnect_0_sdram_s1_address),       //    s1.address
		.az_be_n        (~mm_interconnect_0_sdram_s1_byteenable),   //      .byteenable_n
		.az_cs          (mm_interconnect_0_sdram_s1_chipselect),    //      .chipselect
		.az_data        (mm_interconnect_0_sdram_s1_writedata),     //      .writedata
		.az_rd_n        (~mm_interconnect_0_sdram_s1_read),         //      .read_n
		.az_wr_n        (~mm_interconnect_0_sdram_s1_write),        //      .write_n
		.za_data        (mm_interconnect_0_sdram_s1_readdata),      //      .readdata
		.za_valid       (mm_interconnect_0_sdram_s1_readdatavalid), //      .readdatavalid
		.za_waitrequest (mm_interconnect_0_sdram_s1_waitrequest),   //      .waitrequest
		.zs_addr        (sdram_addr),                               //  wire.export
		.zs_ba          (sdram_ba),                                 //      .export
		.zs_cas_n       (sdram_cas_n),                              //      .export
		.zs_cke         (sdram_cke),                                //      .export
		.zs_cs_n        (sdram_cs_n),                               //      .export
		.zs_dq          (sdram_dq),                                 //      .export
		.zs_dqm         (sdram_dqm),                                //      .export
		.zs_ras_n       (sdram_ras_n),                              //      .export
		.zs_we_n        (sdram_we_n)                                //      .export
	);

	altera_avalon_mm_bridge #(
		.DATA_WIDTH        (16),
		.SYMBOL_WIDTH      (8),
		.ADDRESS_WIDTH     (26),
		.BURSTCOUNT_WIDTH  (10),
		.PIPELINE_COMMAND  (1),
		.PIPELINE_RESPONSE (1)
	) sdram_bridge (
		.clk              (clk_clk),                          //   clk.clk
		.reset            (rst_controller_reset_out_reset),   // reset.reset
		.s0_waitrequest   (sdram_bridge_slave_waitrequest),   //    s0.waitrequest
		.s0_readdata      (sdram_bridge_slave_readdata),      //      .readdata
		.s0_readdatavalid (sdram_bridge_slave_readdatavalid), //      .readdatavalid
		.s0_burstcount    (sdram_bridge_slave_burstcount),    //      .burstcount
		.s0_writedata     (sdram_bridge_slave_writedata),     //      .writedata
		.s0_address       (sdram_bridge_slave_address),       //      .address
		.s0_write         (sdram_bridge_slave_write),         //      .write
		.s0_read          (sdram_bridge_slave_read),          //      .read
		.s0_byteenable    (sdram_bridge_slave_byteenable),    //      .byteenable
		.s0_debugaccess   (sdram_bridge_slave_debugaccess),   //      .debugaccess
		.m0_waitrequest   (sdram_bridge_m0_waitrequest),      //    m0.waitrequest
		.m0_readdata      (sdram_bridge_m0_readdata),         //      .readdata
		.m0_readdatavalid (sdram_bridge_m0_readdatavalid),    //      .readdatavalid
		.m0_burstcount    (sdram_bridge_m0_burstcount),       //      .burstcount
		.m0_writedata     (sdram_bridge_m0_writedata),        //      .writedata
		.m0_address       (sdram_bridge_m0_address),          //      .address
		.m0_write         (sdram_bridge_m0_write),            //      .write
		.m0_read          (sdram_bridge_m0_read),             //      .read
		.m0_byteenable    (sdram_bridge_m0_byteenable),       //      .byteenable
		.m0_debugaccess   (sdram_bridge_m0_debugaccess)       //      .debugaccess
	);

	system_qsys_sysid sysid (
		.clock    (clk_clk),                                        //           clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                //         reset.reset_n
		.readdata (mm_interconnect_0_sysid_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_0_sysid_control_slave_address)   //              .address
	);

	avalon_mm #(
		.width (3)
	) mm_bridge_touch (
		.clk50M           (clk_clk),                                                  //   clock_sink.clk
		.rst_n            (~rst_controller_reset_out_reset),                          //   reset_sink.reset_n
		.avalon_write     (mm_interconnect_0_mm_bridge_touch_avalon_slave_write),     // avalon_slave.write
		.avalon_read      (mm_interconnect_0_mm_bridge_touch_avalon_slave_read),      //             .read
		.avalon_writedata (mm_interconnect_0_mm_bridge_touch_avalon_slave_writedata), //             .writedata
		.avalon_readdata  (mm_interconnect_0_mm_bridge_touch_avalon_slave_readdata),  //             .readdata
		.avalon_address   (mm_interconnect_0_mm_bridge_touch_avalon_slave_address),   //             .address
		.write            (touch_write),                                              //  conduit_end.export
		.read             (touch_read),                                               //             .export
		.writedata        (touch_writedata),                                          //             .export
		.readdata         (touch_readdata),                                           //             .export
		.address          (touch_address)                                             //             .export
	);

	avalon_mm #(
		.width (3)
	) mm_bridge_seg (
		.clk50M           (clk_clk),                                                //   clock_sink.clk
		.rst_n            (~rst_controller_reset_out_reset),                        //   reset_sink.reset_n
		.avalon_write     (mm_interconnect_0_mm_bridge_seg_avalon_slave_write),     // avalon_slave.write
		.avalon_read      (mm_interconnect_0_mm_bridge_seg_avalon_slave_read),      //             .read
		.avalon_writedata (mm_interconnect_0_mm_bridge_seg_avalon_slave_writedata), //             .writedata
		.avalon_readdata  (mm_interconnect_0_mm_bridge_seg_avalon_slave_readdata),  //             .readdata
		.avalon_address   (mm_interconnect_0_mm_bridge_seg_avalon_slave_address),   //             .address
		.write            (seg_write),                                              //  conduit_end.export
		.read             (seg_read),                                               //             .export
		.writedata        (seg_writedata),                                          //             .export
		.readdata         (seg_readdata),                                           //             .export
		.address          (seg_address)                                             //             .export
	);

	avalon_mm #(
		.width (3)
	) mm_bridge_remote (
		.clk50M           (clk_clk),                                                   //   clock_sink.clk
		.rst_n            (~rst_controller_reset_out_reset),                           //   reset_sink.reset_n
		.avalon_write     (mm_interconnect_0_mm_bridge_remote_avalon_slave_write),     // avalon_slave.write
		.avalon_read      (mm_interconnect_0_mm_bridge_remote_avalon_slave_read),      //             .read
		.avalon_writedata (mm_interconnect_0_mm_bridge_remote_avalon_slave_writedata), //             .writedata
		.avalon_readdata  (mm_interconnect_0_mm_bridge_remote_avalon_slave_readdata),  //             .readdata
		.avalon_address   (mm_interconnect_0_mm_bridge_remote_avalon_slave_address),   //             .address
		.write            (remote_write),                                              //  conduit_end.export
		.read             (remote_read),                                               //             .export
		.writedata        (remote_writedata),                                          //             .export
		.readdata         (remote_readdata),                                           //             .export
		.address          (remote_address)                                             //             .export
	);

	avalon_mm #(
		.width (3)
	) mm_bridge_adda (
		.clk50M           (clk_clk),                                                 //   clock_sink.clk
		.rst_n            (~rst_controller_reset_out_reset),                         //   reset_sink.reset_n
		.avalon_write     (mm_interconnect_0_mm_bridge_adda_avalon_slave_write),     // avalon_slave.write
		.avalon_read      (mm_interconnect_0_mm_bridge_adda_avalon_slave_read),      //             .read
		.avalon_writedata (mm_interconnect_0_mm_bridge_adda_avalon_slave_writedata), //             .writedata
		.avalon_readdata  (mm_interconnect_0_mm_bridge_adda_avalon_slave_readdata),  //             .readdata
		.avalon_address   (mm_interconnect_0_mm_bridge_adda_avalon_slave_address),   //             .address
		.write            (adda_write),                                              //  conduit_end.export
		.read             (adda_read),                                               //             .export
		.writedata        (adda_writedata),                                          //             .export
		.readdata         (adda_readdata),                                           //             .export
		.address          (adda_address)                                             //             .export
	);

	system_qsys_pio_touch_int pio_touch_int (
		.clk        (clk_clk),                                       //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),               //               reset.reset_n
		.address    (mm_interconnect_0_pio_touch_int_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_pio_touch_int_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_pio_touch_int_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_pio_touch_int_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_pio_touch_int_s1_readdata),   //                    .readdata
		.in_port    (touch_int_export),                              // external_connection.export
		.irq        (irq_mapper_receiver3_irq)                       //                 irq.irq
	);

	system_qsys_pio_back pio_back (
		.clk        (clk_clk),                                  //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),          //               reset.reset_n
		.address    (mm_interconnect_0_pio_back_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_pio_back_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_pio_back_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_pio_back_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_pio_back_s1_readdata),   //                    .readdata
		.in_port    (back_export),                              // external_connection.export
		.irq        (irq_mapper_receiver4_irq)                  //                 irq.irq
	);

	system_qsys_pio_key pio_key (
		.clk      (clk_clk),                               //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),       //               reset.reset_n
		.address  (mm_interconnect_0_pio_key_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_pio_key_s1_readdata), //                    .readdata
		.in_port  (key_export)                             // external_connection.export
	);

	system_qsys_pio_led pio_led (
		.clk        (clk_clk),                                 //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_0_pio_led_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_pio_led_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_pio_led_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_pio_led_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_pio_led_s1_readdata),   //                    .readdata
		.out_port   (led_export)                               // external_connection.export
	);

	system_qsys_pio_buzzer pio_buzzer (
		.clk        (clk_clk),                                    //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),            //               reset.reset_n
		.address    (mm_interconnect_0_pio_buzzer_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_pio_buzzer_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_pio_buzzer_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_pio_buzzer_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_pio_buzzer_s1_readdata),   //                    .readdata
		.out_port   (buzzer_export)                               // external_connection.export
	);

	system_qsys_uart uart (
		.clk           (clk_clk),                                 //                 clk.clk
		.reset_n       (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address       (mm_interconnect_0_uart_s1_address),       //                  s1.address
		.begintransfer (mm_interconnect_0_uart_s1_begintransfer), //                    .begintransfer
		.chipselect    (mm_interconnect_0_uart_s1_chipselect),    //                    .chipselect
		.read_n        (~mm_interconnect_0_uart_s1_read),         //                    .read_n
		.write_n       (~mm_interconnect_0_uart_s1_write),        //                    .write_n
		.writedata     (mm_interconnect_0_uart_s1_writedata),     //                    .writedata
		.readdata      (mm_interconnect_0_uart_s1_readdata),      //                    .readdata
		.dataavailable (),                                        //                    .dataavailable
		.readyfordata  (),                                        //                    .readyfordata
		.rxd           (uart_rxd),                                // external_connection.export
		.txd           (uart_txd),                                //                    .export
		.irq           (irq_mapper_receiver2_irq)                 //                 irq.irq
	);

	system_qsys_pio_buzzer i2c_scl (
		.clk        (clk_clk),                                 //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_0_i2c_scl_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_i2c_scl_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_i2c_scl_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_i2c_scl_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_i2c_scl_s1_readdata),   //                    .readdata
		.out_port   (i2c_scl_export)                           // external_connection.export
	);

	system_qsys_i2c_sda i2c_sda (
		.clk        (clk_clk),                                 //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_0_i2c_sda_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_i2c_sda_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_i2c_sda_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_i2c_sda_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_i2c_sda_s1_readdata),   //                    .readdata
		.bidir_port (i2c_sda_export)                           // external_connection.export
	);

	system_qsys_pio_paint pio_paint (
		.clk        (clk_clk),                                   //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),           //               reset.reset_n
		.address    (mm_interconnect_0_pio_paint_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_pio_paint_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_pio_paint_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_pio_paint_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_pio_paint_s1_readdata),   //                    .readdata
		.in_port    (paint_export),                              // external_connection.export
		.irq        (irq_mapper_receiver5_irq)                   //                 irq.irq
	);

	system_qsys_pio_buzzer pio_ov5640_en (
		.clk        (clk_clk),                                       //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),               //               reset.reset_n
		.address    (mm_interconnect_0_pio_ov5640_en_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_pio_ov5640_en_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_pio_ov5640_en_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_pio_ov5640_en_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_pio_ov5640_en_s1_readdata),   //                    .readdata
		.out_port   (ov5640_en_export)                               // external_connection.export
	);

	system_qsys_pio_ov5640_id pio_ov5640_id (
		.clk      (clk_clk),                                     //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),             //               reset.reset_n
		.address  (mm_interconnect_0_pio_ov5640_id_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_pio_ov5640_id_s1_readdata), //                    .readdata
		.in_port  (ov5640_id_export)                             // external_connection.export
	);

	system_qsys_alt_vip_cl_scl_0 #(
		.SYMBOLS_IN_SEQ      (1),
		.SYMBOLS_IN_PAR      (3),
		.BITS_PER_SYMBOL     (8),
		.EXTRA_PIPELINING    (0),
		.IS_422              (0),
		.NO_BLANKING         (1),
		.MAX_IN_WIDTH        (800),
		.MAX_IN_HEIGHT       (480),
		.MAX_OUT_WIDTH       (1280),
		.MAX_OUT_HEIGHT      (800),
		.RUNTIME_CONTROL     (1),
		.ALWAYS_DOWNSCALE    (0),
		.ALGORITHM_NAME      ("NEAREST_NEIGHBOUR"),
		.DEFAULT_EDGE_THRESH (7),
		.DEFAULT_UPPER_BLUR  (15),
		.DEFAULT_LOWER_BLUR  (0),
		.ENABLE_FIR          (0),
		.ARE_IDENTICAL       (0),
		.V_TAPS              (8),
		.V_PHASES            (16),
		.H_TAPS              (8),
		.H_PHASES            (16),
		.V_SIGNED            (1),
		.V_INTEGER_BITS      (1),
		.V_FRACTION_BITS     (7),
		.H_SIGNED            (1),
		.H_INTEGER_BITS      (1),
		.H_FRACTION_BITS     (7),
		.PRESERVE_BITS       (0),
		.LOAD_AT_RUNTIME     (0),
		.V_BANKS             (1),
		.V_SYMMETRIC         (0),
		.V_FUNCTION          ("LANCZOS_2"),
		.V_COEFF_FILE        ("<enter file name (including full path)>"),
		.H_BANKS             (1),
		.H_SYMMETRIC         (0),
		.H_FUNCTION          ("LANCZOS_2"),
		.H_COEFF_FILE        ("<enter file name (including full path)>"),
		.IS_420              (0)
	) alt_vip_cl_scl_0 (
		.main_clock            (clk_clk),                                                  // main_clock.clk
		.main_reset            (rst_controller_reset_out_reset),                           // main_reset.reset
		.din_data              (vip_scl_din_data),                                         //        din.data
		.din_valid             (vip_scl_din_valid),                                        //           .valid
		.din_startofpacket     (vip_scl_din_startofpacket),                                //           .startofpacket
		.din_endofpacket       (vip_scl_din_endofpacket),                                  //           .endofpacket
		.din_ready             (vip_scl_din_ready),                                        //           .ready
		.dout_data             (vip_scl_dout_data),                                        //       dout.data
		.dout_valid            (vip_scl_dout_valid),                                       //           .valid
		.dout_startofpacket    (vip_scl_dout_startofpacket),                               //           .startofpacket
		.dout_endofpacket      (vip_scl_dout_endofpacket),                                 //           .endofpacket
		.dout_ready            (vip_scl_dout_ready),                                       //           .ready
		.control_address       (mm_interconnect_0_alt_vip_cl_scl_0_control_address),       //    control.address
		.control_byteenable    (mm_interconnect_0_alt_vip_cl_scl_0_control_byteenable),    //           .byteenable
		.control_write         (mm_interconnect_0_alt_vip_cl_scl_0_control_write),         //           .write
		.control_writedata     (mm_interconnect_0_alt_vip_cl_scl_0_control_writedata),     //           .writedata
		.control_read          (mm_interconnect_0_alt_vip_cl_scl_0_control_read),          //           .read
		.control_readdata      (mm_interconnect_0_alt_vip_cl_scl_0_control_readdata),      //           .readdata
		.control_readdatavalid (mm_interconnect_0_alt_vip_cl_scl_0_control_readdatavalid), //           .readdatavalid
		.control_waitrequest   (mm_interconnect_0_alt_vip_cl_scl_0_control_waitrequest)    //           .waitrequest
	);

	system_qsys_pio_buzzer pio_mlcd_cs_n (
		.clk        (clk_clk),                                       //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),               //               reset.reset_n
		.address    (mm_interconnect_0_pio_mlcd_cs_n_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_pio_mlcd_cs_n_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_pio_mlcd_cs_n_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_pio_mlcd_cs_n_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_pio_mlcd_cs_n_s1_readdata),   //                    .readdata
		.out_port   (mlcd_cs_n_export)                               // external_connection.export
	);

	system_qsys_pio_buzzer pio_mlcd_wr_n (
		.clk        (clk_clk),                                       //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),               //               reset.reset_n
		.address    (mm_interconnect_0_pio_mlcd_wr_n_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_pio_mlcd_wr_n_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_pio_mlcd_wr_n_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_pio_mlcd_wr_n_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_pio_mlcd_wr_n_s1_readdata),   //                    .readdata
		.out_port   (mlcd_wr_n_export)                               // external_connection.export
	);

	system_qsys_pio_buzzer pio_mlcd_rd_n (
		.clk        (clk_clk),                                       //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),               //               reset.reset_n
		.address    (mm_interconnect_0_pio_mlcd_rd_n_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_pio_mlcd_rd_n_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_pio_mlcd_rd_n_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_pio_mlcd_rd_n_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_pio_mlcd_rd_n_s1_readdata),   //                    .readdata
		.out_port   (mlcd_rd_n_export)                               // external_connection.export
	);

	system_qsys_pio_buzzer pio_mlcd_rst_n (
		.clk        (clk_clk),                                        //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                //               reset.reset_n
		.address    (mm_interconnect_0_pio_mlcd_rst_n_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_pio_mlcd_rst_n_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_pio_mlcd_rst_n_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_pio_mlcd_rst_n_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_pio_mlcd_rst_n_s1_readdata),   //                    .readdata
		.out_port   (mlcd_rst_n_export)                               // external_connection.export
	);

	system_qsys_pio_buzzer pio_mlcd_rs (
		.clk        (clk_clk),                                     //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),             //               reset.reset_n
		.address    (mm_interconnect_0_pio_mlcd_rs_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_pio_mlcd_rs_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_pio_mlcd_rs_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_pio_mlcd_rs_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_pio_mlcd_rs_s1_readdata),   //                    .readdata
		.out_port   (mlcd_rs_export)                               // external_connection.export
	);

	system_qsys_pio_buzzer pio_mlcd_bl (
		.clk        (clk_clk),                                     //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),             //               reset.reset_n
		.address    (mm_interconnect_0_pio_mlcd_bl_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_pio_mlcd_bl_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_pio_mlcd_bl_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_pio_mlcd_bl_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_pio_mlcd_bl_s1_readdata),   //                    .readdata
		.out_port   (mlcd_bl_export)                               // external_connection.export
	);

	system_qsys_pio_lcd_data_in pio_lcd_data_in (
		.clk      (clk_clk),                                       //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),               //               reset.reset_n
		.address  (mm_interconnect_0_pio_lcd_data_in_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_pio_lcd_data_in_s1_readdata), //                    .readdata
		.in_port  (lcd_data_in_export)                             // external_connection.export
	);

	system_qsys_pio_lcd_data_out pio_lcd_data_out (
		.clk        (clk_clk),                                          //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                  //               reset.reset_n
		.address    (mm_interconnect_0_pio_lcd_data_out_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_pio_lcd_data_out_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_pio_lcd_data_out_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_pio_lcd_data_out_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_pio_lcd_data_out_s1_readdata),   //                    .readdata
		.out_port   (lcd_data_out_export)                               // external_connection.export
	);

	system_qsys_pio_buzzer pio_lcd_data_dir (
		.clk        (clk_clk),                                          //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                  //               reset.reset_n
		.address    (mm_interconnect_0_pio_lcd_data_dir_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_pio_lcd_data_dir_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_pio_lcd_data_dir_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_pio_lcd_data_dir_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_pio_lcd_data_dir_s1_readdata),   //                    .readdata
		.out_port   (lcd_data_dir_export)                               // external_connection.export
	);

	system_qsys_pio_buzzer pio_lcd_init_done (
		.clk        (clk_clk),                                           //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                   //               reset.reset_n
		.address    (mm_interconnect_0_pio_lcd_init_done_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_pio_lcd_init_done_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_pio_lcd_init_done_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_pio_lcd_init_done_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_pio_lcd_init_done_s1_readdata),   //                    .readdata
		.out_port   (lcd_init_done_export)                               // external_connection.export
	);

	system_qsys_pio_lcd_data_out pio_lcd_id (
		.clk        (clk_clk),                                    //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),            //               reset.reset_n
		.address    (mm_interconnect_0_pio_lcd_id_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_pio_lcd_id_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_pio_lcd_id_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_pio_lcd_id_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_pio_lcd_id_s1_readdata),   //                    .readdata
		.out_port   (lcd_id_export)                               // external_connection.export
	);

	system_qsys_pio_buzzer pio_mdc (
		.clk        (clk_clk),                                 //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_0_pio_mdc_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_pio_mdc_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_pio_mdc_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_pio_mdc_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_pio_mdc_s1_readdata),   //                    .readdata
		.out_port   (eth_mdc_export)                           // external_connection.export
	);

	system_qsys_i2c_sda pio_mdio (
		.clk        (clk_clk),                                  //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),          //               reset.reset_n
		.address    (mm_interconnect_0_pio_mdio_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_pio_mdio_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_pio_mdio_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_pio_mdio_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_pio_mdio_s1_readdata),   //                    .readdata
		.bidir_port (eth_mdio_export)                           // external_connection.export
	);

	system_qsys_pio_sd_cs pio_sd_cs (
		.clk        (clk_clk),                                   //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),           //               reset.reset_n
		.address    (mm_interconnect_0_pio_sd_cs_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_pio_sd_cs_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_pio_sd_cs_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_pio_sd_cs_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_pio_sd_cs_s1_readdata),   //                    .readdata
		.out_port   (sd_cs_export)                               // external_connection.export
	);

	system_qsys_pio_sd_cs pio_sd_clk (
		.clk        (clk_clk),                                    //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),            //               reset.reset_n
		.address    (mm_interconnect_0_pio_sd_clk_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_pio_sd_clk_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_pio_sd_clk_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_pio_sd_clk_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_pio_sd_clk_s1_readdata),   //                    .readdata
		.out_port   (sd_clk_export)                               // external_connection.export
	);

	system_qsys_pio_sd_cs pio_sd_mosi (
		.clk        (clk_clk),                                     //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),             //               reset.reset_n
		.address    (mm_interconnect_0_pio_sd_mosi_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_pio_sd_mosi_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_pio_sd_mosi_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_pio_sd_mosi_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_pio_sd_mosi_s1_readdata),   //                    .readdata
		.out_port   (sd_mosi_export)                               // external_connection.export
	);

	system_qsys_pio_ov5640_id pio_sd_miso (
		.clk      (clk_clk),                                   //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),           //               reset.reset_n
		.address  (mm_interconnect_0_pio_sd_miso_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_pio_sd_miso_s1_readdata), //                    .readdata
		.in_port  (sd_miso_export)                             // external_connection.export
	);

	system_qsys_pio_buzzer pio_page_paint_flag (
		.clk        (clk_clk),                                             //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                     //               reset.reset_n
		.address    (mm_interconnect_0_pio_page_paint_flag_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_pio_page_paint_flag_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_pio_page_paint_flag_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_pio_page_paint_flag_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_pio_page_paint_flag_s1_readdata),   //                    .readdata
		.out_port   (page_paint_flag_export)                               // external_connection.export
	);

	system_qsys_pio_buzzer pio_audio_sel (
		.clk        (clk_clk),                                       //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),               //               reset.reset_n
		.address    (mm_interconnect_0_pio_audio_sel_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_pio_audio_sel_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_pio_audio_sel_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_pio_audio_sel_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_pio_audio_sel_s1_readdata),   //                    .readdata
		.out_port   (audio_sel_export)                               // external_connection.export
	);

	system_qsys_mm_interconnect_0 mm_interconnect_0 (
		.clk_clk_clk                               (clk_clk),                                                   //                             clk_clk.clk
		.nios2_reset_n_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                            // nios2_reset_n_reset_bridge_in_reset.reset
		.nios2_data_master_address                 (nios2_data_master_address),                                 //                   nios2_data_master.address
		.nios2_data_master_waitrequest             (nios2_data_master_waitrequest),                             //                                    .waitrequest
		.nios2_data_master_byteenable              (nios2_data_master_byteenable),                              //                                    .byteenable
		.nios2_data_master_read                    (nios2_data_master_read),                                    //                                    .read
		.nios2_data_master_readdata                (nios2_data_master_readdata),                                //                                    .readdata
		.nios2_data_master_readdatavalid           (nios2_data_master_readdatavalid),                           //                                    .readdatavalid
		.nios2_data_master_write                   (nios2_data_master_write),                                   //                                    .write
		.nios2_data_master_writedata               (nios2_data_master_writedata),                               //                                    .writedata
		.nios2_data_master_debugaccess             (nios2_data_master_debugaccess),                             //                                    .debugaccess
		.nios2_instruction_master_address          (nios2_instruction_master_address),                          //            nios2_instruction_master.address
		.nios2_instruction_master_waitrequest      (nios2_instruction_master_waitrequest),                      //                                    .waitrequest
		.nios2_instruction_master_read             (nios2_instruction_master_read),                             //                                    .read
		.nios2_instruction_master_readdata         (nios2_instruction_master_readdata),                         //                                    .readdata
		.nios2_instruction_master_readdatavalid    (nios2_instruction_master_readdatavalid),                    //                                    .readdatavalid
		.sdram_bridge_m0_address                   (sdram_bridge_m0_address),                                   //                     sdram_bridge_m0.address
		.sdram_bridge_m0_waitrequest               (sdram_bridge_m0_waitrequest),                               //                                    .waitrequest
		.sdram_bridge_m0_burstcount                (sdram_bridge_m0_burstcount),                                //                                    .burstcount
		.sdram_bridge_m0_byteenable                (sdram_bridge_m0_byteenable),                                //                                    .byteenable
		.sdram_bridge_m0_read                      (sdram_bridge_m0_read),                                      //                                    .read
		.sdram_bridge_m0_readdata                  (sdram_bridge_m0_readdata),                                  //                                    .readdata
		.sdram_bridge_m0_readdatavalid             (sdram_bridge_m0_readdatavalid),                             //                                    .readdatavalid
		.sdram_bridge_m0_write                     (sdram_bridge_m0_write),                                     //                                    .write
		.sdram_bridge_m0_writedata                 (sdram_bridge_m0_writedata),                                 //                                    .writedata
		.sdram_bridge_m0_debugaccess               (sdram_bridge_m0_debugaccess),                               //                                    .debugaccess
		.alt_vip_cl_scl_0_control_address          (mm_interconnect_0_alt_vip_cl_scl_0_control_address),        //            alt_vip_cl_scl_0_control.address
		.alt_vip_cl_scl_0_control_write            (mm_interconnect_0_alt_vip_cl_scl_0_control_write),          //                                    .write
		.alt_vip_cl_scl_0_control_read             (mm_interconnect_0_alt_vip_cl_scl_0_control_read),           //                                    .read
		.alt_vip_cl_scl_0_control_readdata         (mm_interconnect_0_alt_vip_cl_scl_0_control_readdata),       //                                    .readdata
		.alt_vip_cl_scl_0_control_writedata        (mm_interconnect_0_alt_vip_cl_scl_0_control_writedata),      //                                    .writedata
		.alt_vip_cl_scl_0_control_byteenable       (mm_interconnect_0_alt_vip_cl_scl_0_control_byteenable),     //                                    .byteenable
		.alt_vip_cl_scl_0_control_readdatavalid    (mm_interconnect_0_alt_vip_cl_scl_0_control_readdatavalid),  //                                    .readdatavalid
		.alt_vip_cl_scl_0_control_waitrequest      (mm_interconnect_0_alt_vip_cl_scl_0_control_waitrequest),    //                                    .waitrequest
		.epcs_flash_epcs_control_port_address      (mm_interconnect_0_epcs_flash_epcs_control_port_address),    //        epcs_flash_epcs_control_port.address
		.epcs_flash_epcs_control_port_write        (mm_interconnect_0_epcs_flash_epcs_control_port_write),      //                                    .write
		.epcs_flash_epcs_control_port_read         (mm_interconnect_0_epcs_flash_epcs_control_port_read),       //                                    .read
		.epcs_flash_epcs_control_port_readdata     (mm_interconnect_0_epcs_flash_epcs_control_port_readdata),   //                                    .readdata
		.epcs_flash_epcs_control_port_writedata    (mm_interconnect_0_epcs_flash_epcs_control_port_writedata),  //                                    .writedata
		.epcs_flash_epcs_control_port_chipselect   (mm_interconnect_0_epcs_flash_epcs_control_port_chipselect), //                                    .chipselect
		.i2c_scl_s1_address                        (mm_interconnect_0_i2c_scl_s1_address),                      //                          i2c_scl_s1.address
		.i2c_scl_s1_write                          (mm_interconnect_0_i2c_scl_s1_write),                        //                                    .write
		.i2c_scl_s1_readdata                       (mm_interconnect_0_i2c_scl_s1_readdata),                     //                                    .readdata
		.i2c_scl_s1_writedata                      (mm_interconnect_0_i2c_scl_s1_writedata),                    //                                    .writedata
		.i2c_scl_s1_chipselect                     (mm_interconnect_0_i2c_scl_s1_chipselect),                   //                                    .chipselect
		.i2c_sda_s1_address                        (mm_interconnect_0_i2c_sda_s1_address),                      //                          i2c_sda_s1.address
		.i2c_sda_s1_write                          (mm_interconnect_0_i2c_sda_s1_write),                        //                                    .write
		.i2c_sda_s1_readdata                       (mm_interconnect_0_i2c_sda_s1_readdata),                     //                                    .readdata
		.i2c_sda_s1_writedata                      (mm_interconnect_0_i2c_sda_s1_writedata),                    //                                    .writedata
		.i2c_sda_s1_chipselect                     (mm_interconnect_0_i2c_sda_s1_chipselect),                   //                                    .chipselect
		.jtag_uart_avalon_jtag_slave_address       (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),     //         jtag_uart_avalon_jtag_slave.address
		.jtag_uart_avalon_jtag_slave_write         (mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),       //                                    .write
		.jtag_uart_avalon_jtag_slave_read          (mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),        //                                    .read
		.jtag_uart_avalon_jtag_slave_readdata      (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),    //                                    .readdata
		.jtag_uart_avalon_jtag_slave_writedata     (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),   //                                    .writedata
		.jtag_uart_avalon_jtag_slave_waitrequest   (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest), //                                    .waitrequest
		.jtag_uart_avalon_jtag_slave_chipselect    (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),  //                                    .chipselect
		.mm_bridge_adda_avalon_slave_address       (mm_interconnect_0_mm_bridge_adda_avalon_slave_address),     //         mm_bridge_adda_avalon_slave.address
		.mm_bridge_adda_avalon_slave_write         (mm_interconnect_0_mm_bridge_adda_avalon_slave_write),       //                                    .write
		.mm_bridge_adda_avalon_slave_read          (mm_interconnect_0_mm_bridge_adda_avalon_slave_read),        //                                    .read
		.mm_bridge_adda_avalon_slave_readdata      (mm_interconnect_0_mm_bridge_adda_avalon_slave_readdata),    //                                    .readdata
		.mm_bridge_adda_avalon_slave_writedata     (mm_interconnect_0_mm_bridge_adda_avalon_slave_writedata),   //                                    .writedata
		.mm_bridge_remote_avalon_slave_address     (mm_interconnect_0_mm_bridge_remote_avalon_slave_address),   //       mm_bridge_remote_avalon_slave.address
		.mm_bridge_remote_avalon_slave_write       (mm_interconnect_0_mm_bridge_remote_avalon_slave_write),     //                                    .write
		.mm_bridge_remote_avalon_slave_read        (mm_interconnect_0_mm_bridge_remote_avalon_slave_read),      //                                    .read
		.mm_bridge_remote_avalon_slave_readdata    (mm_interconnect_0_mm_bridge_remote_avalon_slave_readdata),  //                                    .readdata
		.mm_bridge_remote_avalon_slave_writedata   (mm_interconnect_0_mm_bridge_remote_avalon_slave_writedata), //                                    .writedata
		.mm_bridge_seg_avalon_slave_address        (mm_interconnect_0_mm_bridge_seg_avalon_slave_address),      //          mm_bridge_seg_avalon_slave.address
		.mm_bridge_seg_avalon_slave_write          (mm_interconnect_0_mm_bridge_seg_avalon_slave_write),        //                                    .write
		.mm_bridge_seg_avalon_slave_read           (mm_interconnect_0_mm_bridge_seg_avalon_slave_read),         //                                    .read
		.mm_bridge_seg_avalon_slave_readdata       (mm_interconnect_0_mm_bridge_seg_avalon_slave_readdata),     //                                    .readdata
		.mm_bridge_seg_avalon_slave_writedata      (mm_interconnect_0_mm_bridge_seg_avalon_slave_writedata),    //                                    .writedata
		.mm_bridge_touch_avalon_slave_address      (mm_interconnect_0_mm_bridge_touch_avalon_slave_address),    //        mm_bridge_touch_avalon_slave.address
		.mm_bridge_touch_avalon_slave_write        (mm_interconnect_0_mm_bridge_touch_avalon_slave_write),      //                                    .write
		.mm_bridge_touch_avalon_slave_read         (mm_interconnect_0_mm_bridge_touch_avalon_slave_read),       //                                    .read
		.mm_bridge_touch_avalon_slave_readdata     (mm_interconnect_0_mm_bridge_touch_avalon_slave_readdata),   //                                    .readdata
		.mm_bridge_touch_avalon_slave_writedata    (mm_interconnect_0_mm_bridge_touch_avalon_slave_writedata),  //                                    .writedata
		.nios2_jtag_debug_module_address           (mm_interconnect_0_nios2_jtag_debug_module_address),         //             nios2_jtag_debug_module.address
		.nios2_jtag_debug_module_write             (mm_interconnect_0_nios2_jtag_debug_module_write),           //                                    .write
		.nios2_jtag_debug_module_read              (mm_interconnect_0_nios2_jtag_debug_module_read),            //                                    .read
		.nios2_jtag_debug_module_readdata          (mm_interconnect_0_nios2_jtag_debug_module_readdata),        //                                    .readdata
		.nios2_jtag_debug_module_writedata         (mm_interconnect_0_nios2_jtag_debug_module_writedata),       //                                    .writedata
		.nios2_jtag_debug_module_byteenable        (mm_interconnect_0_nios2_jtag_debug_module_byteenable),      //                                    .byteenable
		.nios2_jtag_debug_module_waitrequest       (mm_interconnect_0_nios2_jtag_debug_module_waitrequest),     //                                    .waitrequest
		.nios2_jtag_debug_module_debugaccess       (mm_interconnect_0_nios2_jtag_debug_module_debugaccess),     //                                    .debugaccess
		.pio_audio_sel_s1_address                  (mm_interconnect_0_pio_audio_sel_s1_address),                //                    pio_audio_sel_s1.address
		.pio_audio_sel_s1_write                    (mm_interconnect_0_pio_audio_sel_s1_write),                  //                                    .write
		.pio_audio_sel_s1_readdata                 (mm_interconnect_0_pio_audio_sel_s1_readdata),               //                                    .readdata
		.pio_audio_sel_s1_writedata                (mm_interconnect_0_pio_audio_sel_s1_writedata),              //                                    .writedata
		.pio_audio_sel_s1_chipselect               (mm_interconnect_0_pio_audio_sel_s1_chipselect),             //                                    .chipselect
		.pio_back_s1_address                       (mm_interconnect_0_pio_back_s1_address),                     //                         pio_back_s1.address
		.pio_back_s1_write                         (mm_interconnect_0_pio_back_s1_write),                       //                                    .write
		.pio_back_s1_readdata                      (mm_interconnect_0_pio_back_s1_readdata),                    //                                    .readdata
		.pio_back_s1_writedata                     (mm_interconnect_0_pio_back_s1_writedata),                   //                                    .writedata
		.pio_back_s1_chipselect                    (mm_interconnect_0_pio_back_s1_chipselect),                  //                                    .chipselect
		.pio_buzzer_s1_address                     (mm_interconnect_0_pio_buzzer_s1_address),                   //                       pio_buzzer_s1.address
		.pio_buzzer_s1_write                       (mm_interconnect_0_pio_buzzer_s1_write),                     //                                    .write
		.pio_buzzer_s1_readdata                    (mm_interconnect_0_pio_buzzer_s1_readdata),                  //                                    .readdata
		.pio_buzzer_s1_writedata                   (mm_interconnect_0_pio_buzzer_s1_writedata),                 //                                    .writedata
		.pio_buzzer_s1_chipselect                  (mm_interconnect_0_pio_buzzer_s1_chipselect),                //                                    .chipselect
		.pio_key_s1_address                        (mm_interconnect_0_pio_key_s1_address),                      //                          pio_key_s1.address
		.pio_key_s1_readdata                       (mm_interconnect_0_pio_key_s1_readdata),                     //                                    .readdata
		.pio_lcd_data_dir_s1_address               (mm_interconnect_0_pio_lcd_data_dir_s1_address),             //                 pio_lcd_data_dir_s1.address
		.pio_lcd_data_dir_s1_write                 (mm_interconnect_0_pio_lcd_data_dir_s1_write),               //                                    .write
		.pio_lcd_data_dir_s1_readdata              (mm_interconnect_0_pio_lcd_data_dir_s1_readdata),            //                                    .readdata
		.pio_lcd_data_dir_s1_writedata             (mm_interconnect_0_pio_lcd_data_dir_s1_writedata),           //                                    .writedata
		.pio_lcd_data_dir_s1_chipselect            (mm_interconnect_0_pio_lcd_data_dir_s1_chipselect),          //                                    .chipselect
		.pio_lcd_data_in_s1_address                (mm_interconnect_0_pio_lcd_data_in_s1_address),              //                  pio_lcd_data_in_s1.address
		.pio_lcd_data_in_s1_readdata               (mm_interconnect_0_pio_lcd_data_in_s1_readdata),             //                                    .readdata
		.pio_lcd_data_out_s1_address               (mm_interconnect_0_pio_lcd_data_out_s1_address),             //                 pio_lcd_data_out_s1.address
		.pio_lcd_data_out_s1_write                 (mm_interconnect_0_pio_lcd_data_out_s1_write),               //                                    .write
		.pio_lcd_data_out_s1_readdata              (mm_interconnect_0_pio_lcd_data_out_s1_readdata),            //                                    .readdata
		.pio_lcd_data_out_s1_writedata             (mm_interconnect_0_pio_lcd_data_out_s1_writedata),           //                                    .writedata
		.pio_lcd_data_out_s1_chipselect            (mm_interconnect_0_pio_lcd_data_out_s1_chipselect),          //                                    .chipselect
		.pio_lcd_id_s1_address                     (mm_interconnect_0_pio_lcd_id_s1_address),                   //                       pio_lcd_id_s1.address
		.pio_lcd_id_s1_write                       (mm_interconnect_0_pio_lcd_id_s1_write),                     //                                    .write
		.pio_lcd_id_s1_readdata                    (mm_interconnect_0_pio_lcd_id_s1_readdata),                  //                                    .readdata
		.pio_lcd_id_s1_writedata                   (mm_interconnect_0_pio_lcd_id_s1_writedata),                 //                                    .writedata
		.pio_lcd_id_s1_chipselect                  (mm_interconnect_0_pio_lcd_id_s1_chipselect),                //                                    .chipselect
		.pio_lcd_init_done_s1_address              (mm_interconnect_0_pio_lcd_init_done_s1_address),            //                pio_lcd_init_done_s1.address
		.pio_lcd_init_done_s1_write                (mm_interconnect_0_pio_lcd_init_done_s1_write),              //                                    .write
		.pio_lcd_init_done_s1_readdata             (mm_interconnect_0_pio_lcd_init_done_s1_readdata),           //                                    .readdata
		.pio_lcd_init_done_s1_writedata            (mm_interconnect_0_pio_lcd_init_done_s1_writedata),          //                                    .writedata
		.pio_lcd_init_done_s1_chipselect           (mm_interconnect_0_pio_lcd_init_done_s1_chipselect),         //                                    .chipselect
		.pio_led_s1_address                        (mm_interconnect_0_pio_led_s1_address),                      //                          pio_led_s1.address
		.pio_led_s1_write                          (mm_interconnect_0_pio_led_s1_write),                        //                                    .write
		.pio_led_s1_readdata                       (mm_interconnect_0_pio_led_s1_readdata),                     //                                    .readdata
		.pio_led_s1_writedata                      (mm_interconnect_0_pio_led_s1_writedata),                    //                                    .writedata
		.pio_led_s1_chipselect                     (mm_interconnect_0_pio_led_s1_chipselect),                   //                                    .chipselect
		.pio_mdc_s1_address                        (mm_interconnect_0_pio_mdc_s1_address),                      //                          pio_mdc_s1.address
		.pio_mdc_s1_write                          (mm_interconnect_0_pio_mdc_s1_write),                        //                                    .write
		.pio_mdc_s1_readdata                       (mm_interconnect_0_pio_mdc_s1_readdata),                     //                                    .readdata
		.pio_mdc_s1_writedata                      (mm_interconnect_0_pio_mdc_s1_writedata),                    //                                    .writedata
		.pio_mdc_s1_chipselect                     (mm_interconnect_0_pio_mdc_s1_chipselect),                   //                                    .chipselect
		.pio_mdio_s1_address                       (mm_interconnect_0_pio_mdio_s1_address),                     //                         pio_mdio_s1.address
		.pio_mdio_s1_write                         (mm_interconnect_0_pio_mdio_s1_write),                       //                                    .write
		.pio_mdio_s1_readdata                      (mm_interconnect_0_pio_mdio_s1_readdata),                    //                                    .readdata
		.pio_mdio_s1_writedata                     (mm_interconnect_0_pio_mdio_s1_writedata),                   //                                    .writedata
		.pio_mdio_s1_chipselect                    (mm_interconnect_0_pio_mdio_s1_chipselect),                  //                                    .chipselect
		.pio_mlcd_bl_s1_address                    (mm_interconnect_0_pio_mlcd_bl_s1_address),                  //                      pio_mlcd_bl_s1.address
		.pio_mlcd_bl_s1_write                      (mm_interconnect_0_pio_mlcd_bl_s1_write),                    //                                    .write
		.pio_mlcd_bl_s1_readdata                   (mm_interconnect_0_pio_mlcd_bl_s1_readdata),                 //                                    .readdata
		.pio_mlcd_bl_s1_writedata                  (mm_interconnect_0_pio_mlcd_bl_s1_writedata),                //                                    .writedata
		.pio_mlcd_bl_s1_chipselect                 (mm_interconnect_0_pio_mlcd_bl_s1_chipselect),               //                                    .chipselect
		.pio_mlcd_cs_n_s1_address                  (mm_interconnect_0_pio_mlcd_cs_n_s1_address),                //                    pio_mlcd_cs_n_s1.address
		.pio_mlcd_cs_n_s1_write                    (mm_interconnect_0_pio_mlcd_cs_n_s1_write),                  //                                    .write
		.pio_mlcd_cs_n_s1_readdata                 (mm_interconnect_0_pio_mlcd_cs_n_s1_readdata),               //                                    .readdata
		.pio_mlcd_cs_n_s1_writedata                (mm_interconnect_0_pio_mlcd_cs_n_s1_writedata),              //                                    .writedata
		.pio_mlcd_cs_n_s1_chipselect               (mm_interconnect_0_pio_mlcd_cs_n_s1_chipselect),             //                                    .chipselect
		.pio_mlcd_rd_n_s1_address                  (mm_interconnect_0_pio_mlcd_rd_n_s1_address),                //                    pio_mlcd_rd_n_s1.address
		.pio_mlcd_rd_n_s1_write                    (mm_interconnect_0_pio_mlcd_rd_n_s1_write),                  //                                    .write
		.pio_mlcd_rd_n_s1_readdata                 (mm_interconnect_0_pio_mlcd_rd_n_s1_readdata),               //                                    .readdata
		.pio_mlcd_rd_n_s1_writedata                (mm_interconnect_0_pio_mlcd_rd_n_s1_writedata),              //                                    .writedata
		.pio_mlcd_rd_n_s1_chipselect               (mm_interconnect_0_pio_mlcd_rd_n_s1_chipselect),             //                                    .chipselect
		.pio_mlcd_rs_s1_address                    (mm_interconnect_0_pio_mlcd_rs_s1_address),                  //                      pio_mlcd_rs_s1.address
		.pio_mlcd_rs_s1_write                      (mm_interconnect_0_pio_mlcd_rs_s1_write),                    //                                    .write
		.pio_mlcd_rs_s1_readdata                   (mm_interconnect_0_pio_mlcd_rs_s1_readdata),                 //                                    .readdata
		.pio_mlcd_rs_s1_writedata                  (mm_interconnect_0_pio_mlcd_rs_s1_writedata),                //                                    .writedata
		.pio_mlcd_rs_s1_chipselect                 (mm_interconnect_0_pio_mlcd_rs_s1_chipselect),               //                                    .chipselect
		.pio_mlcd_rst_n_s1_address                 (mm_interconnect_0_pio_mlcd_rst_n_s1_address),               //                   pio_mlcd_rst_n_s1.address
		.pio_mlcd_rst_n_s1_write                   (mm_interconnect_0_pio_mlcd_rst_n_s1_write),                 //                                    .write
		.pio_mlcd_rst_n_s1_readdata                (mm_interconnect_0_pio_mlcd_rst_n_s1_readdata),              //                                    .readdata
		.pio_mlcd_rst_n_s1_writedata               (mm_interconnect_0_pio_mlcd_rst_n_s1_writedata),             //                                    .writedata
		.pio_mlcd_rst_n_s1_chipselect              (mm_interconnect_0_pio_mlcd_rst_n_s1_chipselect),            //                                    .chipselect
		.pio_mlcd_wr_n_s1_address                  (mm_interconnect_0_pio_mlcd_wr_n_s1_address),                //                    pio_mlcd_wr_n_s1.address
		.pio_mlcd_wr_n_s1_write                    (mm_interconnect_0_pio_mlcd_wr_n_s1_write),                  //                                    .write
		.pio_mlcd_wr_n_s1_readdata                 (mm_interconnect_0_pio_mlcd_wr_n_s1_readdata),               //                                    .readdata
		.pio_mlcd_wr_n_s1_writedata                (mm_interconnect_0_pio_mlcd_wr_n_s1_writedata),              //                                    .writedata
		.pio_mlcd_wr_n_s1_chipselect               (mm_interconnect_0_pio_mlcd_wr_n_s1_chipselect),             //                                    .chipselect
		.pio_ov5640_en_s1_address                  (mm_interconnect_0_pio_ov5640_en_s1_address),                //                    pio_ov5640_en_s1.address
		.pio_ov5640_en_s1_write                    (mm_interconnect_0_pio_ov5640_en_s1_write),                  //                                    .write
		.pio_ov5640_en_s1_readdata                 (mm_interconnect_0_pio_ov5640_en_s1_readdata),               //                                    .readdata
		.pio_ov5640_en_s1_writedata                (mm_interconnect_0_pio_ov5640_en_s1_writedata),              //                                    .writedata
		.pio_ov5640_en_s1_chipselect               (mm_interconnect_0_pio_ov5640_en_s1_chipselect),             //                                    .chipselect
		.pio_ov5640_id_s1_address                  (mm_interconnect_0_pio_ov5640_id_s1_address),                //                    pio_ov5640_id_s1.address
		.pio_ov5640_id_s1_readdata                 (mm_interconnect_0_pio_ov5640_id_s1_readdata),               //                                    .readdata
		.pio_page_paint_flag_s1_address            (mm_interconnect_0_pio_page_paint_flag_s1_address),          //              pio_page_paint_flag_s1.address
		.pio_page_paint_flag_s1_write              (mm_interconnect_0_pio_page_paint_flag_s1_write),            //                                    .write
		.pio_page_paint_flag_s1_readdata           (mm_interconnect_0_pio_page_paint_flag_s1_readdata),         //                                    .readdata
		.pio_page_paint_flag_s1_writedata          (mm_interconnect_0_pio_page_paint_flag_s1_writedata),        //                                    .writedata
		.pio_page_paint_flag_s1_chipselect         (mm_interconnect_0_pio_page_paint_flag_s1_chipselect),       //                                    .chipselect
		.pio_paint_s1_address                      (mm_interconnect_0_pio_paint_s1_address),                    //                        pio_paint_s1.address
		.pio_paint_s1_write                        (mm_interconnect_0_pio_paint_s1_write),                      //                                    .write
		.pio_paint_s1_readdata                     (mm_interconnect_0_pio_paint_s1_readdata),                   //                                    .readdata
		.pio_paint_s1_writedata                    (mm_interconnect_0_pio_paint_s1_writedata),                  //                                    .writedata
		.pio_paint_s1_chipselect                   (mm_interconnect_0_pio_paint_s1_chipselect),                 //                                    .chipselect
		.pio_sd_clk_s1_address                     (mm_interconnect_0_pio_sd_clk_s1_address),                   //                       pio_sd_clk_s1.address
		.pio_sd_clk_s1_write                       (mm_interconnect_0_pio_sd_clk_s1_write),                     //                                    .write
		.pio_sd_clk_s1_readdata                    (mm_interconnect_0_pio_sd_clk_s1_readdata),                  //                                    .readdata
		.pio_sd_clk_s1_writedata                   (mm_interconnect_0_pio_sd_clk_s1_writedata),                 //                                    .writedata
		.pio_sd_clk_s1_chipselect                  (mm_interconnect_0_pio_sd_clk_s1_chipselect),                //                                    .chipselect
		.pio_sd_cs_s1_address                      (mm_interconnect_0_pio_sd_cs_s1_address),                    //                        pio_sd_cs_s1.address
		.pio_sd_cs_s1_write                        (mm_interconnect_0_pio_sd_cs_s1_write),                      //                                    .write
		.pio_sd_cs_s1_readdata                     (mm_interconnect_0_pio_sd_cs_s1_readdata),                   //                                    .readdata
		.pio_sd_cs_s1_writedata                    (mm_interconnect_0_pio_sd_cs_s1_writedata),                  //                                    .writedata
		.pio_sd_cs_s1_chipselect                   (mm_interconnect_0_pio_sd_cs_s1_chipselect),                 //                                    .chipselect
		.pio_sd_miso_s1_address                    (mm_interconnect_0_pio_sd_miso_s1_address),                  //                      pio_sd_miso_s1.address
		.pio_sd_miso_s1_readdata                   (mm_interconnect_0_pio_sd_miso_s1_readdata),                 //                                    .readdata
		.pio_sd_mosi_s1_address                    (mm_interconnect_0_pio_sd_mosi_s1_address),                  //                      pio_sd_mosi_s1.address
		.pio_sd_mosi_s1_write                      (mm_interconnect_0_pio_sd_mosi_s1_write),                    //                                    .write
		.pio_sd_mosi_s1_readdata                   (mm_interconnect_0_pio_sd_mosi_s1_readdata),                 //                                    .readdata
		.pio_sd_mosi_s1_writedata                  (mm_interconnect_0_pio_sd_mosi_s1_writedata),                //                                    .writedata
		.pio_sd_mosi_s1_chipselect                 (mm_interconnect_0_pio_sd_mosi_s1_chipselect),               //                                    .chipselect
		.pio_touch_int_s1_address                  (mm_interconnect_0_pio_touch_int_s1_address),                //                    pio_touch_int_s1.address
		.pio_touch_int_s1_write                    (mm_interconnect_0_pio_touch_int_s1_write),                  //                                    .write
		.pio_touch_int_s1_readdata                 (mm_interconnect_0_pio_touch_int_s1_readdata),               //                                    .readdata
		.pio_touch_int_s1_writedata                (mm_interconnect_0_pio_touch_int_s1_writedata),              //                                    .writedata
		.pio_touch_int_s1_chipselect               (mm_interconnect_0_pio_touch_int_s1_chipselect),             //                                    .chipselect
		.sdram_s1_address                          (mm_interconnect_0_sdram_s1_address),                        //                            sdram_s1.address
		.sdram_s1_write                            (mm_interconnect_0_sdram_s1_write),                          //                                    .write
		.sdram_s1_read                             (mm_interconnect_0_sdram_s1_read),                           //                                    .read
		.sdram_s1_readdata                         (mm_interconnect_0_sdram_s1_readdata),                       //                                    .readdata
		.sdram_s1_writedata                        (mm_interconnect_0_sdram_s1_writedata),                      //                                    .writedata
		.sdram_s1_byteenable                       (mm_interconnect_0_sdram_s1_byteenable),                     //                                    .byteenable
		.sdram_s1_readdatavalid                    (mm_interconnect_0_sdram_s1_readdatavalid),                  //                                    .readdatavalid
		.sdram_s1_waitrequest                      (mm_interconnect_0_sdram_s1_waitrequest),                    //                                    .waitrequest
		.sdram_s1_chipselect                       (mm_interconnect_0_sdram_s1_chipselect),                     //                                    .chipselect
		.sysid_control_slave_address               (mm_interconnect_0_sysid_control_slave_address),             //                 sysid_control_slave.address
		.sysid_control_slave_readdata              (mm_interconnect_0_sysid_control_slave_readdata),            //                                    .readdata
		.uart_s1_address                           (mm_interconnect_0_uart_s1_address),                         //                             uart_s1.address
		.uart_s1_write                             (mm_interconnect_0_uart_s1_write),                           //                                    .write
		.uart_s1_read                              (mm_interconnect_0_uart_s1_read),                            //                                    .read
		.uart_s1_readdata                          (mm_interconnect_0_uart_s1_readdata),                        //                                    .readdata
		.uart_s1_writedata                         (mm_interconnect_0_uart_s1_writedata),                       //                                    .writedata
		.uart_s1_begintransfer                     (mm_interconnect_0_uart_s1_begintransfer),                   //                                    .begintransfer
		.uart_s1_chipselect                        (mm_interconnect_0_uart_s1_chipselect)                       //                                    .chipselect
	);

	system_qsys_irq_mapper irq_mapper (
		.clk           (clk_clk),                        //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),       // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),       // receiver2.irq
		.receiver3_irq (irq_mapper_receiver3_irq),       // receiver3.irq
		.receiver4_irq (irq_mapper_receiver4_irq),       // receiver4.irq
		.receiver5_irq (irq_mapper_receiver5_irq),       // receiver5.irq
		.sender_irq    (nios2_d_irq_irq)                 //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                      // reset_in0.reset
		.reset_in1      (nios2_jtag_debug_module_reset_reset), // reset_in1.reset
		.clk            (clk_clk),                             //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),      // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req),  //          .reset_req
		.reset_req_in0  (1'b0),                                // (terminated)
		.reset_req_in1  (1'b0),                                // (terminated)
		.reset_in2      (1'b0),                                // (terminated)
		.reset_req_in2  (1'b0),                                // (terminated)
		.reset_in3      (1'b0),                                // (terminated)
		.reset_req_in3  (1'b0),                                // (terminated)
		.reset_in4      (1'b0),                                // (terminated)
		.reset_req_in4  (1'b0),                                // (terminated)
		.reset_in5      (1'b0),                                // (terminated)
		.reset_req_in5  (1'b0),                                // (terminated)
		.reset_in6      (1'b0),                                // (terminated)
		.reset_req_in6  (1'b0),                                // (terminated)
		.reset_in7      (1'b0),                                // (terminated)
		.reset_req_in7  (1'b0),                                // (terminated)
		.reset_in8      (1'b0),                                // (terminated)
		.reset_req_in8  (1'b0),                                // (terminated)
		.reset_in9      (1'b0),                                // (terminated)
		.reset_req_in9  (1'b0),                                // (terminated)
		.reset_in10     (1'b0),                                // (terminated)
		.reset_req_in10 (1'b0),                                // (terminated)
		.reset_in11     (1'b0),                                // (terminated)
		.reset_req_in11 (1'b0),                                // (terminated)
		.reset_in12     (1'b0),                                // (terminated)
		.reset_req_in12 (1'b0),                                // (terminated)
		.reset_in13     (1'b0),                                // (terminated)
		.reset_req_in13 (1'b0),                                // (terminated)
		.reset_in14     (1'b0),                                // (terminated)
		.reset_req_in14 (1'b0),                                // (terminated)
		.reset_in15     (1'b0),                                // (terminated)
		.reset_req_in15 (1'b0)                                 // (terminated)
	);

endmodule
