// qsys.v

// Generated using ACDS version 13.1 162 at 2019.01.23.18:52:37

`timescale 1 ps / 1 ps
module qsys (
		input  wire        clk_clk,              //           clk.clk
		input  wire        reset_reset_n,        //         reset.reset_n
		output wire        epcs_flash_dclk,      //    epcs_flash.dclk
		output wire        epcs_flash_sce,       //              .sce
		output wire        epcs_flash_sdo,       //              .sdo
		input  wire        epcs_flash_data0,     //              .data0
		output wire [15:0] lcd_id_export,        //        lcd_id.export
		output wire        lcd_init_done_export, // lcd_init_done.export
		output wire        mlcd_data_dir_export, // mlcd_data_dir.export
		output wire [15:0] mlcd_data_out_export, // mlcd_data_out.export
		input  wire [15:0] mlcd_data_in_export,  //  mlcd_data_in.export
		output wire        mlcd_bl_export,       //       mlcd_bl.export
		output wire        mlcd_rs_export,       //       mlcd_rs.export
		output wire        mlcd_rst_n_export,    //    mlcd_rst_n.export
		output wire        mlcd_rd_n_export,     //     mlcd_rd_n.export
		output wire        mlcd_wr_n_export,     //     mlcd_wr_n.export
		output wire        mlcd_cs_n_export,     //     mlcd_cs_n.export
		output wire [12:0] sdram_addr,           //         sdram.addr
		output wire [1:0]  sdram_ba,             //              .ba
		output wire        sdram_cas_n,          //              .cas_n
		output wire        sdram_cke,            //              .cke
		output wire        sdram_cs_n,           //              .cs_n
		inout  wire [15:0] sdram_dq,             //              .dq
		output wire [1:0]  sdram_dqm,            //              .dqm
		output wire        sdram_ras_n,          //              .ras_n
		output wire        sdram_we_n            //              .we_n
	);

	wire  [31:0] mm_interconnect_0_pio_lcd_init_done_s1_writedata;           // mm_interconnect_0:pio_lcd_init_done_s1_writedata -> pio_lcd_init_done:writedata
	wire   [1:0] mm_interconnect_0_pio_lcd_init_done_s1_address;             // mm_interconnect_0:pio_lcd_init_done_s1_address -> pio_lcd_init_done:address
	wire         mm_interconnect_0_pio_lcd_init_done_s1_chipselect;          // mm_interconnect_0:pio_lcd_init_done_s1_chipselect -> pio_lcd_init_done:chipselect
	wire         mm_interconnect_0_pio_lcd_init_done_s1_write;               // mm_interconnect_0:pio_lcd_init_done_s1_write -> pio_lcd_init_done:write_n
	wire  [31:0] mm_interconnect_0_pio_lcd_init_done_s1_readdata;            // pio_lcd_init_done:readdata -> mm_interconnect_0:pio_lcd_init_done_s1_readdata
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest;  // jtag_uart:av_waitrequest -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_waitrequest
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata;    // mm_interconnect_0:jtag_uart_avalon_jtag_slave_writedata -> jtag_uart:av_writedata
	wire   [0:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_address;      // mm_interconnect_0:jtag_uart_avalon_jtag_slave_address -> jtag_uart:av_address
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect;   // mm_interconnect_0:jtag_uart_avalon_jtag_slave_chipselect -> jtag_uart:av_chipselect
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_write;        // mm_interconnect_0:jtag_uart_avalon_jtag_slave_write -> jtag_uart:av_write_n
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_read;         // mm_interconnect_0:jtag_uart_avalon_jtag_slave_read -> jtag_uart:av_read_n
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata;     // jtag_uart:av_readdata -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_readdata
	wire  [31:0] mm_interconnect_0_pio_mlcd_bl_s1_writedata;                 // mm_interconnect_0:pio_mlcd_bl_s1_writedata -> pio_mlcd_bl:writedata
	wire   [1:0] mm_interconnect_0_pio_mlcd_bl_s1_address;                   // mm_interconnect_0:pio_mlcd_bl_s1_address -> pio_mlcd_bl:address
	wire         mm_interconnect_0_pio_mlcd_bl_s1_chipselect;                // mm_interconnect_0:pio_mlcd_bl_s1_chipselect -> pio_mlcd_bl:chipselect
	wire         mm_interconnect_0_pio_mlcd_bl_s1_write;                     // mm_interconnect_0:pio_mlcd_bl_s1_write -> pio_mlcd_bl:write_n
	wire  [31:0] mm_interconnect_0_pio_mlcd_bl_s1_readdata;                  // pio_mlcd_bl:readdata -> mm_interconnect_0:pio_mlcd_bl_s1_readdata
	wire         mm_interconnect_0_sdram_s1_waitrequest;                     // sdram:za_waitrequest -> mm_interconnect_0:sdram_s1_waitrequest
	wire  [15:0] mm_interconnect_0_sdram_s1_writedata;                       // mm_interconnect_0:sdram_s1_writedata -> sdram:az_data
	wire  [23:0] mm_interconnect_0_sdram_s1_address;                         // mm_interconnect_0:sdram_s1_address -> sdram:az_addr
	wire         mm_interconnect_0_sdram_s1_chipselect;                      // mm_interconnect_0:sdram_s1_chipselect -> sdram:az_cs
	wire         mm_interconnect_0_sdram_s1_write;                           // mm_interconnect_0:sdram_s1_write -> sdram:az_wr_n
	wire         mm_interconnect_0_sdram_s1_read;                            // mm_interconnect_0:sdram_s1_read -> sdram:az_rd_n
	wire  [15:0] mm_interconnect_0_sdram_s1_readdata;                        // sdram:za_data -> mm_interconnect_0:sdram_s1_readdata
	wire         mm_interconnect_0_sdram_s1_readdatavalid;                   // sdram:za_valid -> mm_interconnect_0:sdram_s1_readdatavalid
	wire   [1:0] mm_interconnect_0_sdram_s1_byteenable;                      // mm_interconnect_0:sdram_s1_byteenable -> sdram:az_be_n
	wire  [31:0] mm_interconnect_0_pio_mlcd_rst_n_s1_writedata;              // mm_interconnect_0:pio_mlcd_rst_n_s1_writedata -> pio_mlcd_rst_n:writedata
	wire   [1:0] mm_interconnect_0_pio_mlcd_rst_n_s1_address;                // mm_interconnect_0:pio_mlcd_rst_n_s1_address -> pio_mlcd_rst_n:address
	wire         mm_interconnect_0_pio_mlcd_rst_n_s1_chipselect;             // mm_interconnect_0:pio_mlcd_rst_n_s1_chipselect -> pio_mlcd_rst_n:chipselect
	wire         mm_interconnect_0_pio_mlcd_rst_n_s1_write;                  // mm_interconnect_0:pio_mlcd_rst_n_s1_write -> pio_mlcd_rst_n:write_n
	wire  [31:0] mm_interconnect_0_pio_mlcd_rst_n_s1_readdata;               // pio_mlcd_rst_n:readdata -> mm_interconnect_0:pio_mlcd_rst_n_s1_readdata
	wire  [31:0] mm_interconnect_0_pio_mlcd_rd_n_s1_writedata;               // mm_interconnect_0:pio_mlcd_rd_n_s1_writedata -> pio_mlcd_rd_n:writedata
	wire   [1:0] mm_interconnect_0_pio_mlcd_rd_n_s1_address;                 // mm_interconnect_0:pio_mlcd_rd_n_s1_address -> pio_mlcd_rd_n:address
	wire         mm_interconnect_0_pio_mlcd_rd_n_s1_chipselect;              // mm_interconnect_0:pio_mlcd_rd_n_s1_chipselect -> pio_mlcd_rd_n:chipselect
	wire         mm_interconnect_0_pio_mlcd_rd_n_s1_write;                   // mm_interconnect_0:pio_mlcd_rd_n_s1_write -> pio_mlcd_rd_n:write_n
	wire  [31:0] mm_interconnect_0_pio_mlcd_rd_n_s1_readdata;                // pio_mlcd_rd_n:readdata -> mm_interconnect_0:pio_mlcd_rd_n_s1_readdata
	wire   [1:0] mm_interconnect_0_pio_mlcd_data_in_s1_address;              // mm_interconnect_0:pio_mlcd_data_in_s1_address -> pio_mlcd_data_in:address
	wire  [31:0] mm_interconnect_0_pio_mlcd_data_in_s1_readdata;             // pio_mlcd_data_in:readdata -> mm_interconnect_0:pio_mlcd_data_in_s1_readdata
	wire         nios2_qsys_instruction_master_waitrequest;                  // mm_interconnect_0:nios2_qsys_instruction_master_waitrequest -> nios2_qsys:i_waitrequest
	wire  [26:0] nios2_qsys_instruction_master_address;                      // nios2_qsys:i_address -> mm_interconnect_0:nios2_qsys_instruction_master_address
	wire         nios2_qsys_instruction_master_read;                         // nios2_qsys:i_read -> mm_interconnect_0:nios2_qsys_instruction_master_read
	wire  [31:0] nios2_qsys_instruction_master_readdata;                     // mm_interconnect_0:nios2_qsys_instruction_master_readdata -> nios2_qsys:i_readdata
	wire         nios2_qsys_instruction_master_readdatavalid;                // mm_interconnect_0:nios2_qsys_instruction_master_readdatavalid -> nios2_qsys:i_readdatavalid
	wire  [31:0] mm_interconnect_0_pio_mlcd_rs_s1_writedata;                 // mm_interconnect_0:pio_mlcd_rs_s1_writedata -> pio_mlcd_rs:writedata
	wire   [1:0] mm_interconnect_0_pio_mlcd_rs_s1_address;                   // mm_interconnect_0:pio_mlcd_rs_s1_address -> pio_mlcd_rs:address
	wire         mm_interconnect_0_pio_mlcd_rs_s1_chipselect;                // mm_interconnect_0:pio_mlcd_rs_s1_chipselect -> pio_mlcd_rs:chipselect
	wire         mm_interconnect_0_pio_mlcd_rs_s1_write;                     // mm_interconnect_0:pio_mlcd_rs_s1_write -> pio_mlcd_rs:write_n
	wire  [31:0] mm_interconnect_0_pio_mlcd_rs_s1_readdata;                  // pio_mlcd_rs:readdata -> mm_interconnect_0:pio_mlcd_rs_s1_readdata
	wire  [31:0] mm_interconnect_0_pio_mlcd_data_out_s1_writedata;           // mm_interconnect_0:pio_mlcd_data_out_s1_writedata -> pio_mlcd_data_out:writedata
	wire   [1:0] mm_interconnect_0_pio_mlcd_data_out_s1_address;             // mm_interconnect_0:pio_mlcd_data_out_s1_address -> pio_mlcd_data_out:address
	wire         mm_interconnect_0_pio_mlcd_data_out_s1_chipselect;          // mm_interconnect_0:pio_mlcd_data_out_s1_chipselect -> pio_mlcd_data_out:chipselect
	wire         mm_interconnect_0_pio_mlcd_data_out_s1_write;               // mm_interconnect_0:pio_mlcd_data_out_s1_write -> pio_mlcd_data_out:write_n
	wire  [31:0] mm_interconnect_0_pio_mlcd_data_out_s1_readdata;            // pio_mlcd_data_out:readdata -> mm_interconnect_0:pio_mlcd_data_out_s1_readdata
	wire  [31:0] mm_interconnect_0_pio_mlcd_wr_n_s1_writedata;               // mm_interconnect_0:pio_mlcd_wr_n_s1_writedata -> pio_mlcd_wr_n:writedata
	wire   [1:0] mm_interconnect_0_pio_mlcd_wr_n_s1_address;                 // mm_interconnect_0:pio_mlcd_wr_n_s1_address -> pio_mlcd_wr_n:address
	wire         mm_interconnect_0_pio_mlcd_wr_n_s1_chipselect;              // mm_interconnect_0:pio_mlcd_wr_n_s1_chipselect -> pio_mlcd_wr_n:chipselect
	wire         mm_interconnect_0_pio_mlcd_wr_n_s1_write;                   // mm_interconnect_0:pio_mlcd_wr_n_s1_write -> pio_mlcd_wr_n:write_n
	wire  [31:0] mm_interconnect_0_pio_mlcd_wr_n_s1_readdata;                // pio_mlcd_wr_n:readdata -> mm_interconnect_0:pio_mlcd_wr_n_s1_readdata
	wire         mm_interconnect_0_nios2_qsys_jtag_debug_module_waitrequest; // nios2_qsys:jtag_debug_module_waitrequest -> mm_interconnect_0:nios2_qsys_jtag_debug_module_waitrequest
	wire  [31:0] mm_interconnect_0_nios2_qsys_jtag_debug_module_writedata;   // mm_interconnect_0:nios2_qsys_jtag_debug_module_writedata -> nios2_qsys:jtag_debug_module_writedata
	wire   [8:0] mm_interconnect_0_nios2_qsys_jtag_debug_module_address;     // mm_interconnect_0:nios2_qsys_jtag_debug_module_address -> nios2_qsys:jtag_debug_module_address
	wire         mm_interconnect_0_nios2_qsys_jtag_debug_module_write;       // mm_interconnect_0:nios2_qsys_jtag_debug_module_write -> nios2_qsys:jtag_debug_module_write
	wire         mm_interconnect_0_nios2_qsys_jtag_debug_module_read;        // mm_interconnect_0:nios2_qsys_jtag_debug_module_read -> nios2_qsys:jtag_debug_module_read
	wire  [31:0] mm_interconnect_0_nios2_qsys_jtag_debug_module_readdata;    // nios2_qsys:jtag_debug_module_readdata -> mm_interconnect_0:nios2_qsys_jtag_debug_module_readdata
	wire         mm_interconnect_0_nios2_qsys_jtag_debug_module_debugaccess; // mm_interconnect_0:nios2_qsys_jtag_debug_module_debugaccess -> nios2_qsys:jtag_debug_module_debugaccess
	wire   [3:0] mm_interconnect_0_nios2_qsys_jtag_debug_module_byteenable;  // mm_interconnect_0:nios2_qsys_jtag_debug_module_byteenable -> nios2_qsys:jtag_debug_module_byteenable
	wire  [31:0] mm_interconnect_0_pio_lcd_id_s1_writedata;                  // mm_interconnect_0:pio_lcd_id_s1_writedata -> pio_lcd_id:writedata
	wire   [1:0] mm_interconnect_0_pio_lcd_id_s1_address;                    // mm_interconnect_0:pio_lcd_id_s1_address -> pio_lcd_id:address
	wire         mm_interconnect_0_pio_lcd_id_s1_chipselect;                 // mm_interconnect_0:pio_lcd_id_s1_chipselect -> pio_lcd_id:chipselect
	wire         mm_interconnect_0_pio_lcd_id_s1_write;                      // mm_interconnect_0:pio_lcd_id_s1_write -> pio_lcd_id:write_n
	wire  [31:0] mm_interconnect_0_pio_lcd_id_s1_readdata;                   // pio_lcd_id:readdata -> mm_interconnect_0:pio_lcd_id_s1_readdata
	wire  [31:0] mm_interconnect_0_epcs_flash_epcs_control_port_writedata;   // mm_interconnect_0:epcs_flash_epcs_control_port_writedata -> epcs_flash:writedata
	wire   [8:0] mm_interconnect_0_epcs_flash_epcs_control_port_address;     // mm_interconnect_0:epcs_flash_epcs_control_port_address -> epcs_flash:address
	wire         mm_interconnect_0_epcs_flash_epcs_control_port_chipselect;  // mm_interconnect_0:epcs_flash_epcs_control_port_chipselect -> epcs_flash:chipselect
	wire         mm_interconnect_0_epcs_flash_epcs_control_port_write;       // mm_interconnect_0:epcs_flash_epcs_control_port_write -> epcs_flash:write_n
	wire         mm_interconnect_0_epcs_flash_epcs_control_port_read;        // mm_interconnect_0:epcs_flash_epcs_control_port_read -> epcs_flash:read_n
	wire  [31:0] mm_interconnect_0_epcs_flash_epcs_control_port_readdata;    // epcs_flash:readdata -> mm_interconnect_0:epcs_flash_epcs_control_port_readdata
	wire         nios2_qsys_data_master_waitrequest;                         // mm_interconnect_0:nios2_qsys_data_master_waitrequest -> nios2_qsys:d_waitrequest
	wire  [31:0] nios2_qsys_data_master_writedata;                           // nios2_qsys:d_writedata -> mm_interconnect_0:nios2_qsys_data_master_writedata
	wire  [26:0] nios2_qsys_data_master_address;                             // nios2_qsys:d_address -> mm_interconnect_0:nios2_qsys_data_master_address
	wire         nios2_qsys_data_master_write;                               // nios2_qsys:d_write -> mm_interconnect_0:nios2_qsys_data_master_write
	wire         nios2_qsys_data_master_read;                                // nios2_qsys:d_read -> mm_interconnect_0:nios2_qsys_data_master_read
	wire  [31:0] nios2_qsys_data_master_readdata;                            // mm_interconnect_0:nios2_qsys_data_master_readdata -> nios2_qsys:d_readdata
	wire         nios2_qsys_data_master_debugaccess;                         // nios2_qsys:jtag_debug_module_debugaccess_to_roms -> mm_interconnect_0:nios2_qsys_data_master_debugaccess
	wire         nios2_qsys_data_master_readdatavalid;                       // mm_interconnect_0:nios2_qsys_data_master_readdatavalid -> nios2_qsys:d_readdatavalid
	wire   [3:0] nios2_qsys_data_master_byteenable;                          // nios2_qsys:d_byteenable -> mm_interconnect_0:nios2_qsys_data_master_byteenable
	wire  [31:0] mm_interconnect_0_pio_mlcd_data_dir_s1_writedata;           // mm_interconnect_0:pio_mlcd_data_dir_s1_writedata -> pio_mlcd_data_dir:writedata
	wire   [1:0] mm_interconnect_0_pio_mlcd_data_dir_s1_address;             // mm_interconnect_0:pio_mlcd_data_dir_s1_address -> pio_mlcd_data_dir:address
	wire         mm_interconnect_0_pio_mlcd_data_dir_s1_chipselect;          // mm_interconnect_0:pio_mlcd_data_dir_s1_chipselect -> pio_mlcd_data_dir:chipselect
	wire         mm_interconnect_0_pio_mlcd_data_dir_s1_write;               // mm_interconnect_0:pio_mlcd_data_dir_s1_write -> pio_mlcd_data_dir:write_n
	wire  [31:0] mm_interconnect_0_pio_mlcd_data_dir_s1_readdata;            // pio_mlcd_data_dir:readdata -> mm_interconnect_0:pio_mlcd_data_dir_s1_readdata
	wire  [31:0] mm_interconnect_0_pio_mlcd_cs_n_s1_writedata;               // mm_interconnect_0:pio_mlcd_cs_n_s1_writedata -> pio_mlcd_cs_n:writedata
	wire   [1:0] mm_interconnect_0_pio_mlcd_cs_n_s1_address;                 // mm_interconnect_0:pio_mlcd_cs_n_s1_address -> pio_mlcd_cs_n:address
	wire         mm_interconnect_0_pio_mlcd_cs_n_s1_chipselect;              // mm_interconnect_0:pio_mlcd_cs_n_s1_chipselect -> pio_mlcd_cs_n:chipselect
	wire         mm_interconnect_0_pio_mlcd_cs_n_s1_write;                   // mm_interconnect_0:pio_mlcd_cs_n_s1_write -> pio_mlcd_cs_n:write_n
	wire  [31:0] mm_interconnect_0_pio_mlcd_cs_n_s1_readdata;                // pio_mlcd_cs_n:readdata -> mm_interconnect_0:pio_mlcd_cs_n_s1_readdata
	wire         irq_mapper_receiver0_irq;                                   // jtag_uart:av_irq -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                                   // epcs_flash:irq -> irq_mapper:receiver1_irq
	wire  [31:0] nios2_qsys_d_irq_irq;                                       // irq_mapper:sender_irq -> nios2_qsys:d_irq
	wire         rst_controller_reset_out_reset;                             // rst_controller:reset_out -> [epcs_flash:reset_n, irq_mapper:reset, jtag_uart:rst_n, mm_interconnect_0:nios2_qsys_reset_n_reset_bridge_in_reset_reset, nios2_qsys:reset_n, pio_lcd_id:reset_n, pio_lcd_init_done:reset_n, pio_mlcd_bl:reset_n, pio_mlcd_cs_n:reset_n, pio_mlcd_data_dir:reset_n, pio_mlcd_data_in:reset_n, pio_mlcd_data_out:reset_n, pio_mlcd_rd_n:reset_n, pio_mlcd_rs:reset_n, pio_mlcd_rst_n:reset_n, pio_mlcd_wr_n:reset_n, rst_translator:in_reset, sdram:reset_n]
	wire         rst_controller_reset_out_reset_req;                         // rst_controller:reset_req -> [epcs_flash:reset_req, nios2_qsys:reset_req, rst_translator:reset_req_in]
	wire         nios2_qsys_jtag_debug_module_reset_reset;                   // nios2_qsys:jtag_debug_module_resetrequest -> rst_controller:reset_in1

	qsys_nios2_qsys nios2_qsys (
		.clk                                   (clk_clk),                                                    //                       clk.clk
		.reset_n                               (~rst_controller_reset_out_reset),                            //                   reset_n.reset_n
		.reset_req                             (rst_controller_reset_out_reset_req),                         //                          .reset_req
		.d_address                             (nios2_qsys_data_master_address),                             //               data_master.address
		.d_byteenable                          (nios2_qsys_data_master_byteenable),                          //                          .byteenable
		.d_read                                (nios2_qsys_data_master_read),                                //                          .read
		.d_readdata                            (nios2_qsys_data_master_readdata),                            //                          .readdata
		.d_waitrequest                         (nios2_qsys_data_master_waitrequest),                         //                          .waitrequest
		.d_write                               (nios2_qsys_data_master_write),                               //                          .write
		.d_writedata                           (nios2_qsys_data_master_writedata),                           //                          .writedata
		.d_readdatavalid                       (nios2_qsys_data_master_readdatavalid),                       //                          .readdatavalid
		.jtag_debug_module_debugaccess_to_roms (nios2_qsys_data_master_debugaccess),                         //                          .debugaccess
		.i_address                             (nios2_qsys_instruction_master_address),                      //        instruction_master.address
		.i_read                                (nios2_qsys_instruction_master_read),                         //                          .read
		.i_readdata                            (nios2_qsys_instruction_master_readdata),                     //                          .readdata
		.i_waitrequest                         (nios2_qsys_instruction_master_waitrequest),                  //                          .waitrequest
		.i_readdatavalid                       (nios2_qsys_instruction_master_readdatavalid),                //                          .readdatavalid
		.d_irq                                 (nios2_qsys_d_irq_irq),                                       //                     d_irq.irq
		.jtag_debug_module_resetrequest        (nios2_qsys_jtag_debug_module_reset_reset),                   //   jtag_debug_module_reset.reset
		.jtag_debug_module_address             (mm_interconnect_0_nios2_qsys_jtag_debug_module_address),     //         jtag_debug_module.address
		.jtag_debug_module_byteenable          (mm_interconnect_0_nios2_qsys_jtag_debug_module_byteenable),  //                          .byteenable
		.jtag_debug_module_debugaccess         (mm_interconnect_0_nios2_qsys_jtag_debug_module_debugaccess), //                          .debugaccess
		.jtag_debug_module_read                (mm_interconnect_0_nios2_qsys_jtag_debug_module_read),        //                          .read
		.jtag_debug_module_readdata            (mm_interconnect_0_nios2_qsys_jtag_debug_module_readdata),    //                          .readdata
		.jtag_debug_module_waitrequest         (mm_interconnect_0_nios2_qsys_jtag_debug_module_waitrequest), //                          .waitrequest
		.jtag_debug_module_write               (mm_interconnect_0_nios2_qsys_jtag_debug_module_write),       //                          .write
		.jtag_debug_module_writedata           (mm_interconnect_0_nios2_qsys_jtag_debug_module_writedata),   //                          .writedata
		.no_ci_readra                          ()                                                            // custom_instruction_master.readra
	);

	qsys_jtag_uart jtag_uart (
		.clk            (clk_clk),                                                   //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                           //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver0_irq)                                   //               irq.irq
	);

	qsys_epcs_flash epcs_flash (
		.clk           (clk_clk),                                                   //               clk.clk
		.reset_n       (~rst_controller_reset_out_reset),                           //             reset.reset_n
		.reset_req     (rst_controller_reset_out_reset_req),                        //                  .reset_req
		.address       (mm_interconnect_0_epcs_flash_epcs_control_port_address),    // epcs_control_port.address
		.chipselect    (mm_interconnect_0_epcs_flash_epcs_control_port_chipselect), //                  .chipselect
		.dataavailable (),                                                          //                  .dataavailable
		.endofpacket   (),                                                          //                  .endofpacket
		.read_n        (~mm_interconnect_0_epcs_flash_epcs_control_port_read),      //                  .read_n
		.readdata      (mm_interconnect_0_epcs_flash_epcs_control_port_readdata),   //                  .readdata
		.readyfordata  (),                                                          //                  .readyfordata
		.write_n       (~mm_interconnect_0_epcs_flash_epcs_control_port_write),     //                  .write_n
		.writedata     (mm_interconnect_0_epcs_flash_epcs_control_port_writedata),  //                  .writedata
		.irq           (irq_mapper_receiver1_irq),                                  //               irq.irq
		.dclk          (epcs_flash_dclk),                                           //          external.export
		.sce           (epcs_flash_sce),                                            //                  .export
		.sdo           (epcs_flash_sdo),                                            //                  .export
		.data0         (epcs_flash_data0)                                           //                  .export
	);

	qsys_pio_mlcd_cs_n pio_mlcd_cs_n (
		.clk        (clk_clk),                                       //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),               //               reset.reset_n
		.address    (mm_interconnect_0_pio_mlcd_cs_n_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_pio_mlcd_cs_n_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_pio_mlcd_cs_n_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_pio_mlcd_cs_n_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_pio_mlcd_cs_n_s1_readdata),   //                    .readdata
		.out_port   (mlcd_cs_n_export)                               // external_connection.export
	);

	qsys_pio_mlcd_cs_n pio_mlcd_wr_n (
		.clk        (clk_clk),                                       //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),               //               reset.reset_n
		.address    (mm_interconnect_0_pio_mlcd_wr_n_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_pio_mlcd_wr_n_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_pio_mlcd_wr_n_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_pio_mlcd_wr_n_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_pio_mlcd_wr_n_s1_readdata),   //                    .readdata
		.out_port   (mlcd_wr_n_export)                               // external_connection.export
	);

	qsys_pio_mlcd_cs_n pio_mlcd_rd_n (
		.clk        (clk_clk),                                       //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),               //               reset.reset_n
		.address    (mm_interconnect_0_pio_mlcd_rd_n_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_pio_mlcd_rd_n_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_pio_mlcd_rd_n_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_pio_mlcd_rd_n_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_pio_mlcd_rd_n_s1_readdata),   //                    .readdata
		.out_port   (mlcd_rd_n_export)                               // external_connection.export
	);

	qsys_pio_mlcd_cs_n pio_mlcd_rst_n (
		.clk        (clk_clk),                                        //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                //               reset.reset_n
		.address    (mm_interconnect_0_pio_mlcd_rst_n_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_pio_mlcd_rst_n_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_pio_mlcd_rst_n_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_pio_mlcd_rst_n_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_pio_mlcd_rst_n_s1_readdata),   //                    .readdata
		.out_port   (mlcd_rst_n_export)                               // external_connection.export
	);

	qsys_pio_mlcd_cs_n pio_mlcd_rs (
		.clk        (clk_clk),                                     //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),             //               reset.reset_n
		.address    (mm_interconnect_0_pio_mlcd_rs_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_pio_mlcd_rs_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_pio_mlcd_rs_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_pio_mlcd_rs_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_pio_mlcd_rs_s1_readdata),   //                    .readdata
		.out_port   (mlcd_rs_export)                               // external_connection.export
	);

	qsys_pio_mlcd_cs_n pio_mlcd_bl (
		.clk        (clk_clk),                                     //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),             //               reset.reset_n
		.address    (mm_interconnect_0_pio_mlcd_bl_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_pio_mlcd_bl_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_pio_mlcd_bl_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_pio_mlcd_bl_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_pio_mlcd_bl_s1_readdata),   //                    .readdata
		.out_port   (mlcd_bl_export)                               // external_connection.export
	);

	qsys_pio_mlcd_data_in pio_mlcd_data_in (
		.clk      (clk_clk),                                        //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                //               reset.reset_n
		.address  (mm_interconnect_0_pio_mlcd_data_in_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_pio_mlcd_data_in_s1_readdata), //                    .readdata
		.in_port  (mlcd_data_in_export)                             // external_connection.export
	);

	qsys_pio_mlcd_data_out pio_mlcd_data_out (
		.clk        (clk_clk),                                           //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                   //               reset.reset_n
		.address    (mm_interconnect_0_pio_mlcd_data_out_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_pio_mlcd_data_out_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_pio_mlcd_data_out_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_pio_mlcd_data_out_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_pio_mlcd_data_out_s1_readdata),   //                    .readdata
		.out_port   (mlcd_data_out_export)                               // external_connection.export
	);

	qsys_pio_mlcd_cs_n pio_mlcd_data_dir (
		.clk        (clk_clk),                                           //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                   //               reset.reset_n
		.address    (mm_interconnect_0_pio_mlcd_data_dir_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_pio_mlcd_data_dir_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_pio_mlcd_data_dir_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_pio_mlcd_data_dir_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_pio_mlcd_data_dir_s1_readdata),   //                    .readdata
		.out_port   (mlcd_data_dir_export)                               // external_connection.export
	);

	qsys_pio_mlcd_cs_n pio_lcd_init_done (
		.clk        (clk_clk),                                           //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                   //               reset.reset_n
		.address    (mm_interconnect_0_pio_lcd_init_done_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_pio_lcd_init_done_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_pio_lcd_init_done_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_pio_lcd_init_done_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_pio_lcd_init_done_s1_readdata),   //                    .readdata
		.out_port   (lcd_init_done_export)                               // external_connection.export
	);

	qsys_pio_mlcd_data_out pio_lcd_id (
		.clk        (clk_clk),                                    //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),            //               reset.reset_n
		.address    (mm_interconnect_0_pio_lcd_id_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_pio_lcd_id_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_pio_lcd_id_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_pio_lcd_id_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_pio_lcd_id_s1_readdata),   //                    .readdata
		.out_port   (lcd_id_export)                               // external_connection.export
	);

	qsys_sdram sdram (
		.clk            (clk_clk),                                  //   clk.clk
		.reset_n        (~rst_controller_reset_out_reset),          // reset.reset_n
		.az_addr        (mm_interconnect_0_sdram_s1_address),       //    s1.address
		.az_be_n        (~mm_interconnect_0_sdram_s1_byteenable),   //      .byteenable_n
		.az_cs          (mm_interconnect_0_sdram_s1_chipselect),    //      .chipselect
		.az_data        (mm_interconnect_0_sdram_s1_writedata),     //      .writedata
		.az_rd_n        (~mm_interconnect_0_sdram_s1_read),         //      .read_n
		.az_wr_n        (~mm_interconnect_0_sdram_s1_write),        //      .write_n
		.za_data        (mm_interconnect_0_sdram_s1_readdata),      //      .readdata
		.za_valid       (mm_interconnect_0_sdram_s1_readdatavalid), //      .readdatavalid
		.za_waitrequest (mm_interconnect_0_sdram_s1_waitrequest),   //      .waitrequest
		.zs_addr        (sdram_addr),                               //  wire.export
		.zs_ba          (sdram_ba),                                 //      .export
		.zs_cas_n       (sdram_cas_n),                              //      .export
		.zs_cke         (sdram_cke),                                //      .export
		.zs_cs_n        (sdram_cs_n),                               //      .export
		.zs_dq          (sdram_dq),                                 //      .export
		.zs_dqm         (sdram_dqm),                                //      .export
		.zs_ras_n       (sdram_ras_n),                              //      .export
		.zs_we_n        (sdram_we_n)                                //      .export
	);

	qsys_mm_interconnect_0 mm_interconnect_0 (
		.clk_clk_clk                                    (clk_clk),                                                    //                                  clk_clk.clk
		.nios2_qsys_reset_n_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                             // nios2_qsys_reset_n_reset_bridge_in_reset.reset
		.nios2_qsys_data_master_address                 (nios2_qsys_data_master_address),                             //                   nios2_qsys_data_master.address
		.nios2_qsys_data_master_waitrequest             (nios2_qsys_data_master_waitrequest),                         //                                         .waitrequest
		.nios2_qsys_data_master_byteenable              (nios2_qsys_data_master_byteenable),                          //                                         .byteenable
		.nios2_qsys_data_master_read                    (nios2_qsys_data_master_read),                                //                                         .read
		.nios2_qsys_data_master_readdata                (nios2_qsys_data_master_readdata),                            //                                         .readdata
		.nios2_qsys_data_master_readdatavalid           (nios2_qsys_data_master_readdatavalid),                       //                                         .readdatavalid
		.nios2_qsys_data_master_write                   (nios2_qsys_data_master_write),                               //                                         .write
		.nios2_qsys_data_master_writedata               (nios2_qsys_data_master_writedata),                           //                                         .writedata
		.nios2_qsys_data_master_debugaccess             (nios2_qsys_data_master_debugaccess),                         //                                         .debugaccess
		.nios2_qsys_instruction_master_address          (nios2_qsys_instruction_master_address),                      //            nios2_qsys_instruction_master.address
		.nios2_qsys_instruction_master_waitrequest      (nios2_qsys_instruction_master_waitrequest),                  //                                         .waitrequest
		.nios2_qsys_instruction_master_read             (nios2_qsys_instruction_master_read),                         //                                         .read
		.nios2_qsys_instruction_master_readdata         (nios2_qsys_instruction_master_readdata),                     //                                         .readdata
		.nios2_qsys_instruction_master_readdatavalid    (nios2_qsys_instruction_master_readdatavalid),                //                                         .readdatavalid
		.epcs_flash_epcs_control_port_address           (mm_interconnect_0_epcs_flash_epcs_control_port_address),     //             epcs_flash_epcs_control_port.address
		.epcs_flash_epcs_control_port_write             (mm_interconnect_0_epcs_flash_epcs_control_port_write),       //                                         .write
		.epcs_flash_epcs_control_port_read              (mm_interconnect_0_epcs_flash_epcs_control_port_read),        //                                         .read
		.epcs_flash_epcs_control_port_readdata          (mm_interconnect_0_epcs_flash_epcs_control_port_readdata),    //                                         .readdata
		.epcs_flash_epcs_control_port_writedata         (mm_interconnect_0_epcs_flash_epcs_control_port_writedata),   //                                         .writedata
		.epcs_flash_epcs_control_port_chipselect        (mm_interconnect_0_epcs_flash_epcs_control_port_chipselect),  //                                         .chipselect
		.jtag_uart_avalon_jtag_slave_address            (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),      //              jtag_uart_avalon_jtag_slave.address
		.jtag_uart_avalon_jtag_slave_write              (mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),        //                                         .write
		.jtag_uart_avalon_jtag_slave_read               (mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),         //                                         .read
		.jtag_uart_avalon_jtag_slave_readdata           (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),     //                                         .readdata
		.jtag_uart_avalon_jtag_slave_writedata          (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),    //                                         .writedata
		.jtag_uart_avalon_jtag_slave_waitrequest        (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest),  //                                         .waitrequest
		.jtag_uart_avalon_jtag_slave_chipselect         (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),   //                                         .chipselect
		.nios2_qsys_jtag_debug_module_address           (mm_interconnect_0_nios2_qsys_jtag_debug_module_address),     //             nios2_qsys_jtag_debug_module.address
		.nios2_qsys_jtag_debug_module_write             (mm_interconnect_0_nios2_qsys_jtag_debug_module_write),       //                                         .write
		.nios2_qsys_jtag_debug_module_read              (mm_interconnect_0_nios2_qsys_jtag_debug_module_read),        //                                         .read
		.nios2_qsys_jtag_debug_module_readdata          (mm_interconnect_0_nios2_qsys_jtag_debug_module_readdata),    //                                         .readdata
		.nios2_qsys_jtag_debug_module_writedata         (mm_interconnect_0_nios2_qsys_jtag_debug_module_writedata),   //                                         .writedata
		.nios2_qsys_jtag_debug_module_byteenable        (mm_interconnect_0_nios2_qsys_jtag_debug_module_byteenable),  //                                         .byteenable
		.nios2_qsys_jtag_debug_module_waitrequest       (mm_interconnect_0_nios2_qsys_jtag_debug_module_waitrequest), //                                         .waitrequest
		.nios2_qsys_jtag_debug_module_debugaccess       (mm_interconnect_0_nios2_qsys_jtag_debug_module_debugaccess), //                                         .debugaccess
		.pio_lcd_id_s1_address                          (mm_interconnect_0_pio_lcd_id_s1_address),                    //                            pio_lcd_id_s1.address
		.pio_lcd_id_s1_write                            (mm_interconnect_0_pio_lcd_id_s1_write),                      //                                         .write
		.pio_lcd_id_s1_readdata                         (mm_interconnect_0_pio_lcd_id_s1_readdata),                   //                                         .readdata
		.pio_lcd_id_s1_writedata                        (mm_interconnect_0_pio_lcd_id_s1_writedata),                  //                                         .writedata
		.pio_lcd_id_s1_chipselect                       (mm_interconnect_0_pio_lcd_id_s1_chipselect),                 //                                         .chipselect
		.pio_lcd_init_done_s1_address                   (mm_interconnect_0_pio_lcd_init_done_s1_address),             //                     pio_lcd_init_done_s1.address
		.pio_lcd_init_done_s1_write                     (mm_interconnect_0_pio_lcd_init_done_s1_write),               //                                         .write
		.pio_lcd_init_done_s1_readdata                  (mm_interconnect_0_pio_lcd_init_done_s1_readdata),            //                                         .readdata
		.pio_lcd_init_done_s1_writedata                 (mm_interconnect_0_pio_lcd_init_done_s1_writedata),           //                                         .writedata
		.pio_lcd_init_done_s1_chipselect                (mm_interconnect_0_pio_lcd_init_done_s1_chipselect),          //                                         .chipselect
		.pio_mlcd_bl_s1_address                         (mm_interconnect_0_pio_mlcd_bl_s1_address),                   //                           pio_mlcd_bl_s1.address
		.pio_mlcd_bl_s1_write                           (mm_interconnect_0_pio_mlcd_bl_s1_write),                     //                                         .write
		.pio_mlcd_bl_s1_readdata                        (mm_interconnect_0_pio_mlcd_bl_s1_readdata),                  //                                         .readdata
		.pio_mlcd_bl_s1_writedata                       (mm_interconnect_0_pio_mlcd_bl_s1_writedata),                 //                                         .writedata
		.pio_mlcd_bl_s1_chipselect                      (mm_interconnect_0_pio_mlcd_bl_s1_chipselect),                //                                         .chipselect
		.pio_mlcd_cs_n_s1_address                       (mm_interconnect_0_pio_mlcd_cs_n_s1_address),                 //                         pio_mlcd_cs_n_s1.address
		.pio_mlcd_cs_n_s1_write                         (mm_interconnect_0_pio_mlcd_cs_n_s1_write),                   //                                         .write
		.pio_mlcd_cs_n_s1_readdata                      (mm_interconnect_0_pio_mlcd_cs_n_s1_readdata),                //                                         .readdata
		.pio_mlcd_cs_n_s1_writedata                     (mm_interconnect_0_pio_mlcd_cs_n_s1_writedata),               //                                         .writedata
		.pio_mlcd_cs_n_s1_chipselect                    (mm_interconnect_0_pio_mlcd_cs_n_s1_chipselect),              //                                         .chipselect
		.pio_mlcd_data_dir_s1_address                   (mm_interconnect_0_pio_mlcd_data_dir_s1_address),             //                     pio_mlcd_data_dir_s1.address
		.pio_mlcd_data_dir_s1_write                     (mm_interconnect_0_pio_mlcd_data_dir_s1_write),               //                                         .write
		.pio_mlcd_data_dir_s1_readdata                  (mm_interconnect_0_pio_mlcd_data_dir_s1_readdata),            //                                         .readdata
		.pio_mlcd_data_dir_s1_writedata                 (mm_interconnect_0_pio_mlcd_data_dir_s1_writedata),           //                                         .writedata
		.pio_mlcd_data_dir_s1_chipselect                (mm_interconnect_0_pio_mlcd_data_dir_s1_chipselect),          //                                         .chipselect
		.pio_mlcd_data_in_s1_address                    (mm_interconnect_0_pio_mlcd_data_in_s1_address),              //                      pio_mlcd_data_in_s1.address
		.pio_mlcd_data_in_s1_readdata                   (mm_interconnect_0_pio_mlcd_data_in_s1_readdata),             //                                         .readdata
		.pio_mlcd_data_out_s1_address                   (mm_interconnect_0_pio_mlcd_data_out_s1_address),             //                     pio_mlcd_data_out_s1.address
		.pio_mlcd_data_out_s1_write                     (mm_interconnect_0_pio_mlcd_data_out_s1_write),               //                                         .write
		.pio_mlcd_data_out_s1_readdata                  (mm_interconnect_0_pio_mlcd_data_out_s1_readdata),            //                                         .readdata
		.pio_mlcd_data_out_s1_writedata                 (mm_interconnect_0_pio_mlcd_data_out_s1_writedata),           //                                         .writedata
		.pio_mlcd_data_out_s1_chipselect                (mm_interconnect_0_pio_mlcd_data_out_s1_chipselect),          //                                         .chipselect
		.pio_mlcd_rd_n_s1_address                       (mm_interconnect_0_pio_mlcd_rd_n_s1_address),                 //                         pio_mlcd_rd_n_s1.address
		.pio_mlcd_rd_n_s1_write                         (mm_interconnect_0_pio_mlcd_rd_n_s1_write),                   //                                         .write
		.pio_mlcd_rd_n_s1_readdata                      (mm_interconnect_0_pio_mlcd_rd_n_s1_readdata),                //                                         .readdata
		.pio_mlcd_rd_n_s1_writedata                     (mm_interconnect_0_pio_mlcd_rd_n_s1_writedata),               //                                         .writedata
		.pio_mlcd_rd_n_s1_chipselect                    (mm_interconnect_0_pio_mlcd_rd_n_s1_chipselect),              //                                         .chipselect
		.pio_mlcd_rs_s1_address                         (mm_interconnect_0_pio_mlcd_rs_s1_address),                   //                           pio_mlcd_rs_s1.address
		.pio_mlcd_rs_s1_write                           (mm_interconnect_0_pio_mlcd_rs_s1_write),                     //                                         .write
		.pio_mlcd_rs_s1_readdata                        (mm_interconnect_0_pio_mlcd_rs_s1_readdata),                  //                                         .readdata
		.pio_mlcd_rs_s1_writedata                       (mm_interconnect_0_pio_mlcd_rs_s1_writedata),                 //                                         .writedata
		.pio_mlcd_rs_s1_chipselect                      (mm_interconnect_0_pio_mlcd_rs_s1_chipselect),                //                                         .chipselect
		.pio_mlcd_rst_n_s1_address                      (mm_interconnect_0_pio_mlcd_rst_n_s1_address),                //                        pio_mlcd_rst_n_s1.address
		.pio_mlcd_rst_n_s1_write                        (mm_interconnect_0_pio_mlcd_rst_n_s1_write),                  //                                         .write
		.pio_mlcd_rst_n_s1_readdata                     (mm_interconnect_0_pio_mlcd_rst_n_s1_readdata),               //                                         .readdata
		.pio_mlcd_rst_n_s1_writedata                    (mm_interconnect_0_pio_mlcd_rst_n_s1_writedata),              //                                         .writedata
		.pio_mlcd_rst_n_s1_chipselect                   (mm_interconnect_0_pio_mlcd_rst_n_s1_chipselect),             //                                         .chipselect
		.pio_mlcd_wr_n_s1_address                       (mm_interconnect_0_pio_mlcd_wr_n_s1_address),                 //                         pio_mlcd_wr_n_s1.address
		.pio_mlcd_wr_n_s1_write                         (mm_interconnect_0_pio_mlcd_wr_n_s1_write),                   //                                         .write
		.pio_mlcd_wr_n_s1_readdata                      (mm_interconnect_0_pio_mlcd_wr_n_s1_readdata),                //                                         .readdata
		.pio_mlcd_wr_n_s1_writedata                     (mm_interconnect_0_pio_mlcd_wr_n_s1_writedata),               //                                         .writedata
		.pio_mlcd_wr_n_s1_chipselect                    (mm_interconnect_0_pio_mlcd_wr_n_s1_chipselect),              //                                         .chipselect
		.sdram_s1_address                               (mm_interconnect_0_sdram_s1_address),                         //                                 sdram_s1.address
		.sdram_s1_write                                 (mm_interconnect_0_sdram_s1_write),                           //                                         .write
		.sdram_s1_read                                  (mm_interconnect_0_sdram_s1_read),                            //                                         .read
		.sdram_s1_readdata                              (mm_interconnect_0_sdram_s1_readdata),                        //                                         .readdata
		.sdram_s1_writedata                             (mm_interconnect_0_sdram_s1_writedata),                       //                                         .writedata
		.sdram_s1_byteenable                            (mm_interconnect_0_sdram_s1_byteenable),                      //                                         .byteenable
		.sdram_s1_readdatavalid                         (mm_interconnect_0_sdram_s1_readdatavalid),                   //                                         .readdatavalid
		.sdram_s1_waitrequest                           (mm_interconnect_0_sdram_s1_waitrequest),                     //                                         .waitrequest
		.sdram_s1_chipselect                            (mm_interconnect_0_sdram_s1_chipselect)                       //                                         .chipselect
	);

	qsys_irq_mapper irq_mapper (
		.clk           (clk_clk),                        //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),       // receiver1.irq
		.sender_irq    (nios2_qsys_d_irq_irq)            //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                           // reset_in0.reset
		.reset_in1      (nios2_qsys_jtag_debug_module_reset_reset), // reset_in1.reset
		.clk            (clk_clk),                                  //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),           // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req),       //          .reset_req
		.reset_req_in0  (1'b0),                                     // (terminated)
		.reset_req_in1  (1'b0),                                     // (terminated)
		.reset_in2      (1'b0),                                     // (terminated)
		.reset_req_in2  (1'b0),                                     // (terminated)
		.reset_in3      (1'b0),                                     // (terminated)
		.reset_req_in3  (1'b0),                                     // (terminated)
		.reset_in4      (1'b0),                                     // (terminated)
		.reset_req_in4  (1'b0),                                     // (terminated)
		.reset_in5      (1'b0),                                     // (terminated)
		.reset_req_in5  (1'b0),                                     // (terminated)
		.reset_in6      (1'b0),                                     // (terminated)
		.reset_req_in6  (1'b0),                                     // (terminated)
		.reset_in7      (1'b0),                                     // (terminated)
		.reset_req_in7  (1'b0),                                     // (terminated)
		.reset_in8      (1'b0),                                     // (terminated)
		.reset_req_in8  (1'b0),                                     // (terminated)
		.reset_in9      (1'b0),                                     // (terminated)
		.reset_req_in9  (1'b0),                                     // (terminated)
		.reset_in10     (1'b0),                                     // (terminated)
		.reset_req_in10 (1'b0),                                     // (terminated)
		.reset_in11     (1'b0),                                     // (terminated)
		.reset_req_in11 (1'b0),                                     // (terminated)
		.reset_in12     (1'b0),                                     // (terminated)
		.reset_req_in12 (1'b0),                                     // (terminated)
		.reset_in13     (1'b0),                                     // (terminated)
		.reset_req_in13 (1'b0),                                     // (terminated)
		.reset_in14     (1'b0),                                     // (terminated)
		.reset_req_in14 (1'b0),                                     // (terminated)
		.reset_in15     (1'b0),                                     // (terminated)
		.reset_req_in15 (1'b0)                                      // (terminated)
	);

endmodule
